`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nBlnHi3Kp5ztG6vZNdMONLkWpVVpg2r7ZP2rdZEfioM4XUkRew1oDSrAozd60ivTx8PLiOPPRAJo
pOZd0llK5g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Kcs1MQe5BgqnN7tbrZMcEiZZSCl175bCFWu5jwqWj4RFDG/n9GjuiwAuZ9v2vQZcAxVE3h5w+TBc
Bk1lc9zc7T3tnbm4qpXepckPAqiTqMURQNO28XRRz5BSiTktDkY/dUGVSA0qxTdPGlkYZSpuFpl6
PjievZtLxEtp4cSEwJE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aG1w9h5Ae0N98iRQuCMUHQUwBA2KqP2Fbb/SCJOtosbKahOePVIWiIrkhbLMsr1/omYs/Q6fEj2G
uYHIEBLZLRANmjJt9kQu/jIzWAf0nK3OJkUCAMefyflw5y403PkpWIAHXqlArlaCVW2gWxzVxt9G
js0j3l7Y2dpahAMg2LgLgWyMj2rS0kjr+fbTwgci9As5Ndo6CDyXo7EcixOTvkWvqwxJaYFbtcFF
K1j0WC1jYCLSiEJ2ZB5/ODVnSmn3AWSksydgQ3iYMKpYPNlAwFN7t7HacZ95HxO8MGoNyjnDje35
EzrNZrAA4vUP8Y6En1JgkF6RLt8PJJfLc+wq+g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BYWKn+AL7Gth8aEXuzL+rpOrNP6Ug8Hc9TpmOLZLrPZ4boPFPd89qpRHOY6mfox3M09mZK4TuSx+
5DykxgtH7Gu2DHCqtg3Tg7eFTAzurR/EqXoPhuHQIzs5Y1T/5WlIb0c4l9CNWdc5TBVfbmKR+x4N
A259tw/6q69OtmAqFiB+p9GY8lyjNDWu07DJlxI2l6wSRYy8YqD7K1OrLRXxY6gaTqDWDXlcO+ia
T5/harPHjTiNAFO8U6YTfRQtNJUrOnNfSAnAtjrlegYGNcEl6u4sqYE/X/Pajk2n+1+KvJ6PR8L9
bdrCByV81f1z88nc1Twl6LUe54VQdfe5W+EOpQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iJnLIMkUEl7Btn7IVUeqK6xbyk9c7fsISctkfj2c6osS1GvgHXWHkJPpNPHTeIth7zUvkUlYB/Jd
M5kNK3leJJj5TaqOLOh+cyWqEGY64EruHImVJasbLaVn3LUh67wEEMFoKhP9/KjqLsL3oFrKnU4i
JzYtVgZoCfaHBaIyRC6wms7z/YKP2Khya0dzmYHMmbdm9k2rL27fVLJcCEMSO1Dsz2D/qXnCFI8T
NHnM3Fv/xF2jOhtDIDqWGakvXk7l+ddg95MJ+5A578jqVX81M0WJwbHlaIJIG5uwIzTI46+pYw0Z
4sgDMkrl/aXSFYB5PU2L4hhVeq7e6c0dqUOVSw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sdiBszQspScY+UIwuaohSbs1PAZL6bemuOZlFLGklUXNsz7r1265PlclnSy9m0ilIWxY0HJkGEtl
Rs/zfRlF9Ag/CEiBQ4lStxiXa4cbOvNwkp9j1BXCYCAbMsw83x+ZvpyoQTXRfcBBvSAbtpFDJ7ar
qlJbO6erRjpDP373GIY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eUV1ae8Aw6l0UtyVDuKmrMQwdVI8vrJTYSKwNJ+/x3fs7qy5B2fVzNE8tFRcie7NykwBpJV9lQNN
iNNcReVBjS/oh7txKer0RVLuw2jQCeQBSixWXwdIra9CsrIF5V2GUuY3dDh9ofaqsgbKSlDNLzzm
0lHhjAw4Nbk9kwoo5NP9xZYaLPCNo4Qqi0A9Px++Zu3V7DcbPDDDQnNEzgQhcN8ilscDyGVOeiHu
/xJbo1lLkpyrDciztvHYqwj9O/kSyF1PikDg8xEaOx1QQVvaz7r51DlXlPCpqCUyFGEeiIrPCMHf
8rf7t9DpvBEVPF3eaofCDfiW9vWmbfgffwtMYg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261312)
`protect data_block
eq7yPN7bOKZcd+PM+uZpJfnCvYwD18XR0ASzeXiyEG6WHH94SM89K6EKzWPQDFiwTPWoQAEUmLub
2JuJBcFcLN/2XQT2vyhhLAir/iGWAplf43evC82ix5WervrBGkWZM1Bq3napD4CVvj2bslrGQnwY
piVhq1sLBjgWjbQXQUqyt6VLzjOftcZEUgqRii9vyMLExsiNBsMdFAt+KjdQvLxxOrn7xPdYf21+
3KZyZ6d2IywVWqqCHL18IzgpiB7mOQsH/MRYCmBbspXVP++vv6jhd/Revdv176e9gC5qKYxrscnw
g16GsQS4+wFBX6KC236HnLv78wDl4D40yuZ0eaVcny+HdHbYwwjvf3yIWPdjmHnRIkg81BEUtpJw
Y3l60AEAjp9fJ2F25jQydBXJo3xqN9QjIa1GvlzIfU0CxYa/tWvC7lWcEuI/xh1F6jl5vUo8xhTS
oV/66GvEDWCEd7JRhCbO+Hm/e/HipCyN7NkSJJazbpmxM8Y5K50h/Mq8Fp1fQMl92i4CimJsO08x
/VYLjdCe5/S5yL4XuDwIqBrDYEYxw3Ktg8S76oZ4svAysfW6W7tqb5ewqzZfl9cn9vldikvwO0qa
7DknKqW63xwj5KkRQsSeSVkXekCD6yVqMD8iMeejZaA+RbrWFXU/ExROrc7UFg8Si8BtnXojK5ZW
h9B36jf2JNuXREE+8kXjaL27cts+txQpIgEV1VHAvagT5hUjtAZGgzCyrhrkzPnq+SR5GZLgkVZB
UI5r0SSkqqIa5vborQSDRnRCiO3WIZL1+drQC5vxfDo7KmSyYwOiQT9kwwJlJ4GbdHry6U6NUh5q
bwqTSrern1mEgT2rCap9U3Nmph0k/IeOKd9LX7HFrdTXbEtdN70taIjR5muCJm5YfzNNr7v+ae1a
eU85rywK7Qe/hEmSCIIZJ3eSvhN4IY+1ET0t0QSE8IqZVfV9ZlQ6pYcY7JP2s3AjdZS1XMfA0IxB
W6+M23nyf0P2IlcdZ+BlWL5xuapwIMCqRwS9YuaZKtifTklRzH3KcEzYjeClSdvPQ0SvYZ4WG0j+
XWtemANyldT1ojA2vqtcvE3RUrpRlao/1aRXCpAOIUISrcYRv0WO7G7rC8xRw7p4TFcAPtMVyv7b
KSw+/dkmJQ4X1R4rffpHiIZWqXnP8UycPIO0HzInank7G8t5dsIegEDGgzX/cWmKVzwAanMh85jy
+jjMryYdZcMon8fCX5cmEnvL5p8FxEWaw6Ek+nIgWrsSHdltFMSrM0UjdFM3FxHZTkQfaHu/uxxk
qUCE5OKoI2Z9HJ2CVpEqDB4RiU4CtLX9cfqqiO+q6+f7jzzpPsBjhyXNForrjuE1XxiwVzFBmgYL
rRp47h3EAxM7gsgDUPZM0hDwE8BX6A9DyPhNOWYGc5mYWviLRoTVd73oQ/J7YAvbIv56bFr0zdWr
cxpNMefDnGJAfFdebyMs2NWZq3l4TwmGR7r21bQOsZkttWKKNUrX5yS2LxRe/AJNTPV0qnVtWrXS
Vr/IAKNxRKLXgKtuwc+bm4svJZK036BN0Rko5MPeGGWaTtl+Rb2jUehCsWtGIdxorEmuO9ES4Muw
rwfcECcfQNSAMUQpkPzvPdiLDiun+b+OBND3GBG2ei+cjNubmTJWaUuN+Mh7UKGjTyoKoap9YrOp
OZLlodtylwJqmAKptmZyoV//PAwk1hZmLq3Lwn/BF2JXOmVwqbXtRwtI3rvVvx13Jq8EcxOEbPbN
YoQ7ybjZ+a2qWzx6h/LGpYoeL4yUWBzTRqwua/hwY+SVeZb/BTiNhLdBAznal7r51BSxtVdyebHw
fzqaINPCPwDbIDObBam25QMJWoaGsmj1Yt71imEZPE0jicMNSNUo1wNFrbHs0V5MnZ1OEwi/cRMg
Nn7LxQ6UGZK2qdmZu4K3lNf9uFefHYZWtXfjBBsZgX0lb24NRwU4MxZQRBaV15fkj+yRQpdGd3YO
VH6qNCY83bXYymREVdeuxGe/gK+wDTsQQDaISslwhDsSwO52Ma2pBffL1UcId1NbUZkezvxZIh+Z
t+f9QiCc7QF6U9Pwxd7RnA9LFW0f4t0GdHof7Z2u2FjfJmpbsBqE2c90GWsHXqQQ6Gl6U1Fa9Ics
AC3xdBpz+CgYPQbVOC5B8ChWPe8QE7rBfdJW2BAOlH7g9YJXpT/n6oweAQn1vihrQ9JRVk59oG/E
cwCsm+BkmFJsGHxqCNivgFGNi/LWNbwYZ10BwL1nAdhhOHRUEU1lzICN/qTj1KwwENFx0mJOOvYZ
ctLWUhEHXbYKw5rLkT91O738GCwegA3Zo8WxgUVvj71TjILbOt7yl0JvtfsUpR3MtRzfxgrwuDMI
BULFeHM6COQdm1BOCJ0SVpxKBuopW9BxKP4DKgPwX7pHAUJ7/hUcmqcJ+HwKH3e6sdkjDmmM0lpk
xWhA7LwytEHv9J1SCOHafMQA3aWJCTOOOzwPMf1qh1RQtVQHBr91DnJvrFmoViLembuJN9tUZMA2
Ucr3xCWFnItVh/QkquMD/A6v7gkcdfFeZBOebfOsLIzwIs/6honjzsCFQCBUCHqXz8tlbnCr+K0U
7xreeBo85N2jMh8EOJ6qOnNv/ORgmt2uTiTrWUUY27L6XB7FhaN+TwFR+oAKN6fvgXD2luuIgzkd
59auWQ/rHLPZFtM0Q2y2vqtpWadg8m1yBN/E125CPhUoL4rPL1BS5/aRwlgNDugHD2P77sYPPvot
lw6XEu9AzGyAkoJUtwizVRh0IG9GtXluxmtTKqaucvtZnJKP4p+75Ypsl4ltD0hcbk0zdqjVMar5
Er4KC6g2xzQbQ1RfsrcOtIm3Mfx0fFB9WZFEkP4dk78HPQJLwukSTMJbw2nMnhXCus9LeSlJ+wwi
B/z6ol6nu5lAnrpLPZ946YxVglpfquX3VAMiqbZW36xomPdv5WgyagX1Uy24O+hG11dgfFw+Y7fw
Kj68ytuSrvk49rVJM/YfAFl6ItZDikGXddV/UeI2f8lZn4QyNYYezKHWkn7wqKSOiJNiuB/FBLNf
/GhfHPmXGXKlOpl0KN9YSpY+N9yYL0PctVeGy6LaBTFm1FqFls/DuKn2CIqIOceyv9/kShOCSSj2
d0DBMDWwUW7JMl65Z+TgRDorxHqjyhJ4DKGxlQ3zZWrnKeE8CT6lFccMA2z84hr6Mm5cA9i/d8ha
cBMcTtJWy9XjPi2oUcS4L06nM9heTu0POBZ/uNRHPrIUKSmnnDfj6qd4FeMNVQQn0wCc1WNFIkm3
8k4wT3CQQLD9T0DbgyZfcICckjQe/TTd7uyvs87+qlkt6bbWPMha7zX0igkELYPNFyI2KJPQlIY4
ocBwv7SKH9E53zxEyY4Xz8PbvbQAJ9T8OPwybcxUsP9AvbCDOc4BdACljJHh0C2On964EZsdNttl
U1dQxC7PPzaaSa9bIjwyupq/oIiQgHE89yxlFZVtaMA/K8PVqCAWYgdgz8XfvfaX+9k2JgxXFMah
I/aYgegcJbWs5sc6USEPhZg2pBYt/03aMZpGSbsR5FwLjLKrSP4pWZd0n45aWlJdbFgIj9GiahVP
Rxkyvg3JUYnzSF6l95+VqqGQT6Vi3VrgNp5SdC58jx/JHMvpthFHbdbW36TMYyHuAn/t2EmuBvFi
0vIGFSIUJPq9l5h+O7526/qizqIb62cXFmgIDkBltg7T7/eWICJNs000Bh82RYSfCSPdkX1hhOEK
1JLW3LcN8/9u/ED8RCgSr6KMND6QoNYqiaWzBvPC6KCFNR6TRu+czbmFGU1kN4nrHfCIZX0WrPuo
kzBcSI9ImXQQX6aGXyfyW/zdwJZG+I+Z1QPXf6XEQIzpsYZXxPssXJUiGSjtu8VoRnsHbCD+iRPu
gvvo3xnHchEVwMpUmHw3HtkMcHbB+CMW2ZVzcIudgB+MIvT14knPz5dvT256q8CEBz7bwuVaipYw
pWQDfik2krHtaojN7dVFIM4dZtNHfbLUdv/ibbxR5uioi0A1bqe7YwLAA4g1y7+cQV/ODuWS01ET
ZsZMGkSvtf5FnhmptUItmncv67tTXCYHNZxDE9Vyb1BSVBxbq+DdvoBUfWRNuX6aELP7yhfGWDq8
g51/4WwdNLOLJNu4GmvGGe31iXl0CBaan4GqW0ZMCpyP6b9AAS9sBtVUKml/lmaQZpOfgz7LbgTh
5eTCI7u2Fawvg+te5N9TdvGAZR9ZKJkTtCMqsL7mnLewzdXudd2CJQVuIBosHE4CaAz8rgQpLEHi
AF9goVCV9n5rM6QZEbB6CPGzBlsweUL/eYIXrt0/9iA0zffdQ4kKYSGqce+TckME+4VBYBqCzexs
wd29raKd/YusSObRqaPvteC6sO3uKRZIi7e9M6t1tfizX3x15a/79SqFuoR2yqZ4hwWcJBDdQfXT
RzL/lI4Sl8wB59NyZl6Hl5JL9Ej0ZXp7+YvwsKHFQe4KYr+w4/4E/mBeaBIi6pmujW/+CM6v2G2/
+Rfp0VRJxVEodILkwLfwBtEX2WGnj1dVW8s9PEx/nquLKkppUrnriWRjHpZCwpgQEhtWtqTTf8Op
ucy6dTnSqOb9uD/b+TGryAtK5W3cLfxMmgN3ARxJhOvP89rdgX4vJN0DsgcxJsW0VLI/QG2iwAnd
X1TcJ3b3ykwAGTY//UeqeuxMmqQ+pKKi9KZ30jo2Px9D7LtEtacog9eCr+z74C3gfnd+IGhvTkPB
aPr+Q21Sp3ictYE+zbXwFM/ExHJZrJdOdOojX23r1qTBPypjF7ryweL6Y8oLmjBdNQBfcblbLOV2
YJNSu5fplo0zs3985h2I6vk02PiZ+cuGmo+jB1nsTUQfXkNW0049r2KDC2Tcc2Ng7oZ95tJRodiU
PtGEuLVF+2uwZkXZAq8bVKWLT4uOEncg6ANwix+DF9YaA0+JJ1HS1xn906Jg5XHmEmA3l0eBW0Lu
hrKOAgCyr0uwLAcpJXXxABct0W8EoKczNdjdHnUW8lUcHpeYVysH6bVNijtj1YU/0pz6LIVnEySv
0qVVDTlOcfrtTMp8RTKScfqyWRu8NR2c/tjD5L1mBFXx9zh0xi3ZRO9ULxdOFeOchiaspXGK/YyA
bYnYFJ5rsWBT0tEGHBiUVreKgCUv/a7Hd/k8+t2GjpDEIRdpM92h31CnSycD/fZ5j8pkXN9iuVCL
jY4JGFchN5z4KZEvBKPNEFdtUPei6I3dpBIciTSCxywon0rXMaWdDgrBxviW4onLKzdhtFcpxceD
5flDB8jC06j7OFf5kaMe8EbFriIWXx1anmXoQ/KDha3kyoZdKEumztejxP3C/gXX8HBXPOm4nW2h
2O9mHjz89dZN6b5u2Lq6htQ5uXEe3Ae58d2FuDoLVhJwEjQpUIMpjO/GmtXhsf9j3s+hq+frR5Dr
hrK8KRpH7PVRYtidUKpGXLvp34XMuc1+IaDUQf4hWsCBl/az19SeHNjjEx0V3lwN0jP1BAi2hCcB
V25uY3gAP0pqHp9Z+0sYFSNrW5AZfDXBF+E3wH3ukW2dtZFgucu472g4oQd+8rkAIHBpPUR/yur0
JOGgdnYQS38wqaOAYz5TGdnMsU+ZXdiWND6c42AtvyiZKunRQFRhZKdjEFEg71Owo5zhh3rJUO4F
vItTaINagve+wF8dKwwcDOEPd0tgvN3HykdmW91wqzUEypDmqeLtAeFcLIkjhF6YEpoB+/GvCA+S
ubqf8GSvFtWmRituS99DpiZTkjBDIwaIQd4MlLyTItP//WhzDnTVIVu7l1Gi5dh+KOnILA0EHHJI
u9tw4LOja2PoZFt+tZ9qsg0MGNF1W3ItNmhd9Fc57iUCNUV3sX2Qdj3UFtQ4Br+W1gu2U5E9K1qj
uJqSqjVk7cQw6MefiymW97bG2v+pBP0m9ye3VG6u/ezX62q78pePi0vTdjeDslaeOHSFXsm/2htr
bongehp4GcXwxsbmukH9IlXqm0tww+TK77U6mlKJ293sesVO2M0Hv2E/TWl6+3qLDn1o6UWkmdPA
yUzWTh+Fgg0j3jqQ64rcz/8KLasU4TflbXz/6ZcENJjAMfUSPMse+O+rAaSvrdtVvJ4fyF7XQ62W
2zTf3gLKtERL8A6STg20B/TaYoVusJX5N3vJrQDydQo3KKEin02MgUNXsHoMv/RXdDX9RD1M5guC
JbAh5TC4SbRat9hFwLF72nK7VPVfDFMYP/o5eQFYAK4eqksZRYdNI8FXLc/N59YOzBiUzVe1uQEt
NLugaBYFJTpr8p5JILP8/lYEFipkfmhS/wnAOIyC5DZDGNHdUlsZiNZCOECdkj5yUSwy/5WP3sNP
00CPIYw+WR09u5cTCI9D925Xv66I/p2UbhVrmsK6V5FnQCn8MaFC+D5EFdh7oGbDbgtqTTHsvTjY
i6Q60lpEt9I9DxfcO+KjDhMpxuDjyLGXwxD27W9jb4jrP7/yKs5/MwQoED8dVddj8S5YiJ49GTCt
CS0lysXUZbjisQ1CyM/LRGCG5peOkAMzC+Y+QFUKw0mD+cFeWbs3M4V7NhtliMUTwTHXp4S0caUu
WzEvY6vNcTf4hNOWRYyUDIdHJ9/i/b2qmAcCZ8dlkE7+3gW/go4Wo9zVGVgx8u5mhSwojlwmnQR5
ma9//EXIBmFKGJaHu9MP/4xKLytRm0dnhXunRlo/R6iNKAgCLWJP8tk04TH+VW6h41cd9QvswsHS
Nh+/RjJTUDODLwNfOvyvXcoWTFZU2nFC/nUfTihD6P/FQFYRFRHJD8OzhzsyoxPLm538bHhEo9hY
87gJHdPG5nzuauIs/aht5KBmo5k0C0WtQReALwa5tHBHfyayjdugsfI56KqNYXG+L1zCfzc9bJFx
m4L0TqxdfZ4hyMLYnatris8f2Mmm9w9zVLHKAPFauCxdx2DEFdWJC9dWBTP9tb61x6c4/0o4sKXa
vNzalnyYO7CRZAaqzNKDQl3MRiDCEw+ltbRQWQRBl/5fADqv70jeUBh1A6F3WCUqraYzmJEQO+hE
/Ax766SAJll+/JztIymDgm95XL9mwwi+ddzXV0fT2KyUbL/GJ9lutqihFnluTKte/2c/VoSd+YKf
pt961zh5aRetJiYYfmnTqfGc6JS7wtxmGNPWOCTpDVOGr6mJ5E9n/pEJHiWCrS6J2z20aUjpiwWe
zAVmMCEots/fgqaGyYE9Z3o4jsVZyukgDzABMDASxqDn+NnM359Lp7hSY3QXAwxrDkC/WvTKNQiK
VJk9GN6cOzwH7xF6WGrfc5Ct20BsK39PGiCMYT3H9b1g0IEF+eC7IkAckfvtiZjhWZBkDHDZXmNI
LaQdt4nu820exVFiofDhoXLIQAF6/n5pgEiyiToFiWryUYujSd7j8D1oPG76KV7nTSKTZS5+SH+P
n/Q8/RU/IDTucKDV4E4Ln4XaiiXTJXMdkc8zdg4fflV6m8znYgMSRmFJM2TkVVO2Ss46D1+qwI1/
MdwxAoD7BwFweYMtpC+dr9ugyIMm8QpBxB+cWk8yN+0bU9Sr4g8afmS/h5lnWCILYMmhTXQFzejx
NCgjBJLdSPOHR8loBLQYOXCbyu40IoyYykskOs82vXTCy+5hQ+XXJyV47Oam93CD87BCWuo2lR1U
CzXhS/owpGy5QJVWT7vKfAjtFPL5QPOBz3WT6IOvVqY8QEq395bFBWqMgoCXrPgeAZoEndYc9JE2
PrbOHNC/7B0zHXjWeIXRCghzJqitb32qpe0jTlXw2vQBR1PEjf4mVY9brqt5PbuM/MJwUUgMMIIB
Yx4zWTsh88gib+v+DVdo+beoh5Cm70wKkLyRl1sPkt9H2hH/0qaLBaPSBk8fUkYO+jvbCJ431wXl
qxquKFQyDuWp6Z4xD7O0QshlsSMm757q0PZDdNY2q7GondqyXygUkmDueo+iWJc5gFeFGP/X75+M
b00UpKYMLkNYvWsxfxsxTOVQ7/EULZaoMHBoz4QzVUy62f1WwMC6NBStVc5F2dCh2GVDDFXya7cw
5chAdBUpP3WWd8+ddJt0gfPO9GniV3LCAU4p+N+JC+R20Wh1JvABrwvwk+6ZqYq8efW+uuJSi49Z
J9NJcSnbq7E8a5R4yKq7rzIWnxuwY1x7Wj92fnTfYwZCvANQAtD2P/hucbBjSTwNEdQIad+zRfgI
RGLwvTpArqX6ZL18HQo5ZyONl/pLv2MNbk4VbcsiAyHkVlTV4qXRbw2t7Qcsd/JzMhJa+3PCUcdA
fAXXjIsghE2Mwcfrztj9pKZAT+G5yJF08FLIDbfGgsGawDwZiOZCPF0obTUUMIZCEgEK1CzmJ9Ax
gW5N+0+4R+DSwZOfR3Ii92mmgTOXJvv+q1fBSTLKIdmzQ8I8WGPn/UdeZH6JpgyyKZlgaxD/86LS
H8qEuJhF37aa1AlQU+kPgmhLFi/YGx7SX6XL/SM9dH6NcvXPZDcSSJtDTuiFSWzVaTrxfBsMBhdH
9h7ny7haWfIAFaRq0h1ZYw+qAf9akNcxjOUpEtA7G+wl11Z8pVTwrh8M3c+U8VmMUBuX/ubscksU
ahWxYEDZ+uqxfHqhlLZgB0q0Z2zhmPS4H15sJvjJMMBqWpH0WAVx7/t0T0bGxHHPa9WsWuKbsQ/n
bVO436HIGyNglzrYQzeW8oUeSyBi0MvaEuVjYpyK2hIfV52nl3aQs8/A1+8jJMBLn1HX3Nc4dOH5
oUSJu/lSxp9+sfD3FJfdzNamcmzWJ5Y2djiqSyVK9BmQiVOCC8XDIucNi5ToDZUEAwVKiDIxirZQ
OICuT/dpx/k1MHHzawQbC21GTWSZs4Wf4tg3ltLaXnuGfHTj2IyVZiJN4Bvoz33BBcguLvIOpWB2
xUKNcYCXf+IQQUqFGgSx2Sin2XszTjefiNQ9XFgcKdqFT4blYhsmMvB/DIgCE+WuW11Cq0t+Pid7
IfYJ63nuy7FKmcHyUUj2n4I4xkd8YLho1RWLHHtufwgqBuKPiAh38wBw6v0zs3j2P9I+NcIWYGy4
3CEBaGbtliQsHZ3Hmgiou3R0/h2uCzxh3TBXErUh4/ozYk3NA4anSaFqvp1kGSIiOluV/CoYnMbU
5OFETH2vANjIUTTK5H4yj8wLcEvvrS8CDcKuTH4U/UsutmCQBle2dkf5WcpIqJEa1z89nF7ldkWF
5S4LE3tzyAEcIaSbG6JNtWHW33TWpu5qeqfwYHChHcu2400dxKQxef0NQmKNQTJhTrEjhbjNeZXP
F7vZp6ToP6a8xV4SjgZJqGFqgh5HkiNPVRHKdAtsKUIX2FzmzWftXFp0hA8juMZkeY2Jxvo3VIKz
F/ImbGpu2ScoZbrQwn9xWCdq27OAjDtjCGrnlZVFf6v6dhb6xhOdN3IEIOXth3CRg+ZwyF2KK17G
JKPyP5d49JpO45eCOP/2MyYu/otbI0mySJPNk2mRR16OcGhyUx44UYFwwxE/ADpvwoOgPJZh6WIk
0I2aDikmPA3JJyDGialpf5GMaiPABKcuzhTJ52Q7fSRXr+DtrYuUClExVO9Wx5GoN8vzAJJ2m+Dr
P0GoNgHuHC+BC/mWbBNB+r7McWWKUKITEl5xgVEw0Bw9piuB6bMrYPh6iQtd41WoncjS7pQYMi2z
62wA1tNW4d1aiq1BK6PFAmVsWhGHD5TJMvErw7f0YsRwyPFezuLdOAEGlQmV0nRkDRefzaSqGoNY
CxtkKHetPT8086V10zQhK6P9YhEFkLVAUjLPHrn4lH04r8xYACRyXcavAxWMlKgCY+bB+x8kwAOU
RCLbsVBx7IqfkeXkn05mwd/MCv0Gfo6uoiv0aRTlDSAdb0tUOmGTb65zkHLFuuO62Y6hutXanymJ
xx02VHsaiRaMUpJ9ntGthrEiesGXYlpTXnfyrLum/5jSNxqbHpeqLl0/K2bKlkvzIWi2M9JQp/ac
eG2Pw337jjjFMV8VLeeNy5uqSY18CuT+fRW56ZjzHizNlnbD5445R10CQdV9aVatoyezNgsg/JsF
vR54hpOX0Lkp7Om9bsUeZjjwvo7huu9+ku1kFVmnQUstMn18MEXD1DxPbvVUUYOu+7t45CNkOSGu
qq7HqqSddo3lIXPy3wDY8QPFd1GMqo8juVlk9njFP2evMXhGOg5I0bcFlCy6gH38dm82djaqAs6u
G8/3+OtX77LScoPLkYIVRU5Ed3m0+uMZjfeAsRwj+obg+OdfJEf2kN+tXE79jCU2DTbn1/iK7vDp
q7aausNtKz7A+i0D/Xz1vrJZ3K8ttQBaR9yENorqEmyrnApFW+rBpmh0h6ts8O6v8B34g1MiTHw5
WOdZFNW6fnvdZrP7+xo39/cz6UMczci+RNEOL3B4DAcwGQfrrgpoWY+JQcB/Fo/SCeHx0bHtBumc
T6o99ME8tlPd4J1fl+g3cZuMWHTTTR8D5lWc76O59WqUXtSSkhupQJfObpRIl0M4Lw4bVp4AUTd3
5zfu7ranf+RDAlmMe335WLjRP+RXilWxERco6jzBJi/NYn8JAGQGVouNpvAyPWtDrbsbR3WXJYBU
PRrlA5uexIk86frj0q5RKPKmR1bfm4i/7Vwl/QukkxPXyvVf/wVX93o5SmMbF3yxbNuN3gGybX3c
G57elayiDYTCfvzo1S2POvf4+bQtBLf8gUR0le90SryQBgBqeJbJgg8pd03rMYe2XVASr0caSNK/
FjTBpJK9njGer0VFkQKPR+1UrL2MTHD+PXwB9PghwY+60+aVV0E1CdfSetuRsrpqBfH16MtuipPQ
OsuRuviYCp9qfYlF1P3z1riDlqKPq1t2qvdWSVino76EmotjXoE7YW3+/NY2XyooVshyF3VCuRZx
pe8yvL0ywelrsQC+ih7fl2+ympiRISzV1c9SSN5ETvrA5Yf85aR/gq1wnFFkxms/a9PaQ5EO8oIg
HgyWcV8joErd5vrBSGA4fqLTPweu86/AZj3aV3GrbrK47eW65sHiyHqMolJmYk2QKt5r2ejVvbeY
fiysCbH51lWRlkB8vd8w6X3Wrf+oOQg+wZ3CM4247QSInv5PfvImDF82BatKrORBqtZaVcH6PSDM
gg3H4vY8Yx83MtALRjM57W3T4nFMiQElnqQeC05ojG/GyiaGlKUzN/87t6sx+1goRBRsb9SgdKvO
5QXC6W99Ru9MY2A6AkCAXRfHYiFktX21SguCTp0HQ1Ef7hgHUFJ079LPluDZO5DBWgQz+OrDQusd
Dle4ZUlkcPx4ACfnk/j+peXLnk0sfaXNuBbue+uGl7A10N4Bf7qQ5/9PTJdWUSxGiEcCOhq6vDCT
mwra8W9FB9OUfk7DfhDQybLtz24r8rgLcEov0ytaD4RHb27h8amknzH+5ptDV1MAVbaHtRsgsn+L
AVT0q4DINdW0WMER/sv+WVU9Z6FBtfbttVTnr3Fh3xAeBS/fCCJV9COWqL13cDEbvNV8EyuzJIO7
u6HJ1mY0knSxR66Olqn9DOi4iyVIREBixjcM/62WfNtWMngsJmSfQ7VSUDGXm7FKR5BlJFAxyXFZ
40is6VfWGnNgrgID1VInxB9cijqyYoIy7AK3BHvOWMi29DICrsXwSWY69h8Xb7uMR7pja09ee7q6
vfVrCE8oCgLkkfjgKmxLw1PeYXJIDZ0FSF4wE30lxyuXISJLokVRndxjSP/v+l/Fh//vkwajMCIn
Qx5kyPD5YjSwAG1e4M8qJ6xWgkDbIJTbd4TmeXUWN9lNeNMAWx+rF6r2fllTjm8hZQydz4Om9ROJ
os6Xl4s5a1ETc/U5pXRkGkA3eTOZWWz2l3z578k8biyjGqROT//ojp6Cys/1XvzHxS8MWlFQvnLc
uaNIFioM1/wDA1wd+YHEbVVuCbiI7m/sCbXkjMGKcVObWHoEJnU3F4lCmlnJDcuN0MhwqbDOUSm6
oD83ZFtLI/QgrcNRMij6WZi3D5cWESFNEpo5yvsEfcBFJfYmhZqPx2bj/md+EwPVILjTlY5MIdVr
YNMuVIHBfFrSuI0cP6d2aT40QnTlhJ6PPQS3opPQeTd7HIK3zPz/wx+VIdlzUKvzB566EMasjeeu
uonCIPrS7zSHzWDx1wJM1EuHI2v7Di5/LsGMHNlL8+nPrrAndEaBbCfLC42fvxnSs1nBoC5p9g6D
zDZrHnskUNDCudCAA/LPPIwBNHOjhnl9N3/PzUgF6lspF04t9uGQIaSFmVtDXM/hgS31CKaxW5N8
jCbw6QIGv40FUG2NeV8NQ4Zu+9RGxbtBLiMN3XNq+sG5VrJxjXBzqPwQdBtS5pD6/kxrmtW0RZMk
wZlufLLy3WaY0ASBf3TleHbBhLwi2F81Hn2MGqWge+V7OTpLljb6bmdQGYbB3zqHs1tF1A0CdZHh
eVi+Yk1v/RTlAUAZigGaXTTr2mVlbVGKfrkbztSmvLx864m5r3Dlg9XGS0j0ctCjaJzEeV7qwEKQ
Cp+fzBso8IJ+WGHsxMAspSqgPya0NT/Um7brym0rMxMuBwKC5OYP4aJKVFWk0Goulm4gs6EVl8k1
AhPuj1HD0kE2sCcEMJrrZY8GgQ30SawF7H0+3d3hMN1B3BO4Eec3/CcD2MpJcWPM58MEfv5mAeE8
WLlMZ4gnJEZntUweD3vYnTbicpHG/lNa3m8gCkfjIUI3xcnBtxMgQA/sxkIJTL/DW2irsgwjuO9o
KE6Tmjqonhy2c2cInm6rwq1wkszOUQ0RhJLUsq+k+rCoPp0EDTP/i9woEjQ9OoSGBUtgxAIVhJ85
OsEBl7j1J8ScFy3DWS5+bMPeBRZwmv8S28ve2lhBZAJOgrRMpHh9q7ANrZJirfCYgTyZrlIONUcG
KiDHVMfyCP0xP47zDwT1Bv4cOMWkNhNWGeqv3sD9I69GFKoDQWiESxuk+7Pk17VAmQEb9FwZng2Z
T92Tpb/T1WDkbU3K86XP7jyP0Yq2O69xeKqWBkpq+LEMjuooKle5k7L2KOm0xY3g/GgYZAjzWOQd
v5s28ou1Vdya5TTs7yHiEOqRm2kaUcSZk7pedmCvh7WsWpNdkRUwq3X1gJCEdOCCm43eaA2nb1O5
GLcHOisUrLHqDGOzyb6wRpYSeHSWufiOkLzLlbt22ALvPZ09uMZdXRWjeSLbrOdClvpfW3sazZ7l
vYiy/Jv81Fx8CX6n8BbuRgq7nilzFbd3KUITqnSsV2F1DNSkjKG3e4CNCEgK1D9eKNfsHW6r3ZyF
Lgb/aWCR6i8zppMad5K67i7WldGAL4BLKwA7wbRPE0p960Ajobq9WrJGVfa9hUxoJtVpVIF+ePbo
SA06PAvZxu3yNhRPNiyPcmlveepnl9bebMivO5WDYg/H8+9WxIk6N954b2lvbTfzyaLeB8z+Lirs
4ydnuOyI6o1pabSLigjAUkaYLkDeATMkIQ7TyyJ1wmRVHttW/OqXKlrNaULcv4tl7WGwJ+1TYaJy
c3cHkZv+J65RehFJRh7RkwJrvTan8jDi+4UkcOAlzI0YCWiJJwvf/MGzP6tvItvaTaJeZsGQDM/6
wVGYcCG8b6+jJ8K76czua81c0NudUP7QkyfF3YgCAdL2GDpkZX0LcfuJD11IwHVT3Xn2n4nV2jOA
0JMjC4B4My3qcb5Y85uejdswee0dRTcpG0yXcMSB3wddt+pLj6No2SJKqaqqRVC35gZs6wp/v7e9
hFod9vf81rFvAbvaEjAeSCywkF6Mhto6k5iRr1bUWjuFNhdVXyQm6Yi5O7du31tY3o8kBHxpfZyn
2BlXso544Gdl1VMVMKzjqvMhbFUeYPbmwiiq5DjSwQSsbKKG4ssHWY7K6iEZzVFgNUKYe8QnmPs7
fB6J4RDF0WY91mOBxuv29meIrpzZz2VrYn8RYYYM95n/PCxk6G0qhpTiSGAph2z07UGsSNcqvdpA
X8lCQHbP3G5pJ2yHjG3rwOu7JQk1NHnrHVP/tW2pHPkn5bYo8sYwl1vHOnOq7DCkV0MJ7xrbiUsZ
D4Kfqmu8juKqpI0eyDbU1YdOem22dlcTu9AhnmchDdwsV4Rz7n6AC2qYirOi+CIXWDiTeWlyqBFQ
tAs2cpujDnrlJjWtARLBOa6HhtgpiG3Om8/Ozd4gU8WQi0WFQaMvJ5oUl/pJ77231nBnRBjbCF8q
d2cs5w3yrB2Lrr5kZT3dvbZ32GVae70P+Zi+VqpCXKqTvQ3HAW+91y9x+aVzUN36rA17B0NbiypY
Iu+3vc7rbUO2pDNKAVnfSlk57IOkG/1133PrrZObpi+3rGgiOc9LGG9zgBx3uBMaz4a8taKHIhWf
Y6cuG48dF2chUfX8JOcP1QVTMTunJJcO61QgPVLm4r1x0TY0/LlF8W2RQKuMZZOnrXS7Vkh3zM9q
ggbDtBNyOVPjjivSZ2f9Rtuf1NgxTO2dAd8LOhgh7FU8Sb7+raEOrlHuwiobmXvOvKZdv/BE79mu
oZxRXQp0pdsdcs/Hv0BgnqLhMM99VkAtPjvtFF/umWTdez1us3dihTYW8EICP9aCjsH1uhSBX86O
gZT7j4MNCHHnM3/2Mrjqmu+9gQ99PAYb+BZm5K2U/lOSOtzQYKf1V6iktgCqX4BSKlo7/J6ezVfp
ZD0kDVw1hP4GWcsUcAtDgOJZpoDw1wSffpF8ImycqjWnSEJGs6HZARQgpwMlwhrk5WbnnYR2lZyc
tx1JSQP7EV61Xh1vMkkPDIiGv3/ufQL6c4/n20pKkbI1kn7eZVnDztH86bhGKovbUeA0Jpr5k4fM
76jT0R2arAhryyFatsuFFsxnqoizKKj9hQnHfn0i1ZQCdiWsmCEo4aR7ZRvjQJbkJJ+5NPK9jQnB
uOReGnquM9ZHjv6jFKP4lcrq4ih0CZ4A+htPaQEVlHHuRkmC2BzjOwFacIdK5jdhrKDpj9wH2WvJ
i3sJdQSfqiyOxYQ4kfxcb7SjQt3rimWfzchuHbmpjSQ+LQqzh3okzt3gqhUaqW0/SO4QZ2c8Kd0h
+JKgFK0DVnOjs5l4K7cN1z1WVxSun89b4zFmqqQX2y7IRYDyAasGKfXKzqdkcYDis7baWMjistc+
X7l4B3OlKiSkXuqRsl9yLZs1c3unainHQ5xO7GhD58XCLg32WsVJNBztssQd69ezE33Idm1V07Z3
NS38mVp5lVJyBJohuNDw/KwxNdqEDTHfbRY8rMspyy9dye94GKmQCK26DTour9ThyyKhjO2gqgCi
qNb68NSx6bw1Qj87LpOkwb+ns7IoiXYRW2kHbO536FXN18Ha0r1M8dhzBq5jnMh35PzK9vMOoKT0
Su2XYQGIhB9It17o7KYSI/vNOi9JwuIfqoPqi7Q8346F/2GQZOJsotYDwpMLlQMAIPtduEvVD0Tw
dZE1N7DHLhy6IzB9BIyoW7jvrkXB1rJBba4EGlVeexiM2NrFDAE5G9ymRO0iaMMV9LJIoTxgR8iu
rCkM+5fM5qJu2I0iuAoHtOzqgvVPei5aAdNeHxqy2UCG5aFdsjz1XB5zV1zxa+KIxYig4EjlgZPW
VRJwgOJpo2myJNQG2411+lODODQDCJjzT48EPGJUqSo79eFp52l4gWutkvAjT66hvoZAlxgeLDyb
RGA2aHetANuDWH1u4fu69V7pyu774f+6Xr+h68sIzrK+4+OGNcP4gi3gFpK6GrGEWSK1gytfqcGR
A7G4coQD5mZmRaxBV3gcJFufAZq17vm0bFiseRhA9dBM2TYgvT/BXBmlhJ7Z+4gaBXNYIG2w36QL
GkXOnhkk5jkjP0/Z62acnki7oADn6Y1Az6peEzQWSy8DFgGdD0GBEvdQzh98uy8MsXmj9OJr1c2a
2aITxs/tIOkItNW6OoD3gJwZmrZ2v594y0hTWvJ4uOHfoDE1TW9BrWgE++hXo07AsR5I6ZflEnaY
/iJjo7Uk2BZUH5EhAmhurPzcQz229f4ngNU6+EpURGVI0Nq1vPkoAy8V9LugMFvLJ+Ku4h0z4xtU
cPiPcjpvNsxVu7fpI84URDKxTPUn9/lO1AadG/sCCMi02jPgoI93ho9tDoThOMuK83xvwI+8Yrcq
H9D1h/95EJmMTo37NDIxOahGQaJaq4XbCJAEXSruilzCUIdWwQmkyGY7pyTiUljLR/hTz2WjA+bQ
fcnJVbZbKTGeyZupT/HfK9g23uQ5ygIuSWjlSt0+Y1V8JAnCg4n3Fc6tFyJGjey6951BeLeJUz1w
L/r3eJO44F7ZJSnOYgQtb+Zx6o/xF6AlSeAdsDiBI58PtKUR0qX7XwvWM/CW90DJpspkw8XRgUko
tqmaKLataY4/lrIgLB8dFLLaVtuqyx9NuURSWolvCWfVw8AT4rhQUPf3LGhbCNi6PDnOV8QJwIZd
IR7/sXq1z7mlKs4smQfpK883Bksyi3OnxVZ3UpSDUJRYdxHv1fhbEs6YOZzNDV/5GMicGLZ+OY+L
Co3U9hkJ4tUCrnt+uOLuZCJDo+Aj8Tin+TPthVF3FQFoQSn37bcBkGmO8PhAxCIkPzD2WfyeI1Hu
ydjASW/PUTQiP5V/6snyv7bN63iq7Jo1k8p6XjweK5TSt3C+rf5JqCg2xBun9XEboqcV5ONnkTGs
4YQ2SLhE7IW2dPwo57Bk+OhqQKhOVSLZ9F3CGzqf3nOIB3RrzK/UxqeYIXc+8V1J+wb7qgf6cf0E
HK1WdZqo+nP2XTYa3Wn61MnIybHaSASmfZxLxxa+brGYKkiCrvUNdPscGBtc1mEvnwBSQQS9F38u
Ckimli5GWreJQkgOyHtRLEhnbVPDP+PLgJFejqV/+2wRaZE2zgja26D6sQEoz0YXD335IGlgx7UL
zRamAxlrHVhDBm6x/Vv42eOOuUHQoTL9umfKLAKqFhBQv8PlZK+5h24OJjtrI/BHqdIsf1pCBbwm
SD7CprtXofbDpIa7ElBdTNvYtQG/xoQD/+bX5P4VOKi7uHJedtCLGCAmybpHzptdU7ltpt9i/CNY
wex0CLkiyoAPO2JexbirEbpyHuYogCtgSgyk5U1Bc8K4qonqBK2MpzgOARfdZRPAFB208N11bl8q
TSgd+srjzcW4Aek6boDRqlPk6Qy7++FMHeOYM64LDQ9r+ASYYSN6OEo1JrgBEgIw46KEh+cT0Aas
FywxeSIsxp1vka1AEnj6YbQUL1H+4cWtZO5VU0BIwtpdlpjpf6461OE1sZyFzE8j63azrdhYWw/6
H8i07DXfF/gXMK/iDNSgge1QP21tmxChT1/EgATQ5LoXbahMyKdq8jSblVXn3HIDakyWWA5w7Z/t
BmfV0m94QQi1JsxBFSKvNwKM0GreSOzXSCMc3OeSaj3piAl+7UDFmAwFK8Samr10/d892upfi5YP
oSxif4ujS5+3LLO2bpvEtrWpBMJlom694wVYxd+0bt9IcSQU6B4XBi0Bt+/gnKiqF+YoQBmJp9sL
3bChxNpegn7GlLdWahv/NUcwpKAQgLC/HjZ+P+XmKDxwGzeyNe3LB6Oboe6t88mdjbVPMK2Iu6tK
fQq5i9eqiKg2bHyNDUW6hiSY8sOBo/6cYKTE1lbmGb5pF0r4m+0uEtwwg9F6+44do9E9h8ieYZ1X
yTk40JFyKR3RMbbD9oCVHydg9S4Hy4ZY7mOpu2GeE84AR+v/8PWfUHmjmVHpihfokQasunmCslOP
Au045WYUSDGZ6QKOoT/YK3COnSdoM7jDcw/TAIP4EzZZ3KzGsuwXFRtF4wAUSfpjL2qfZmkH7+IK
WF0f3GangsNSdEkKtDVm4dibOhXsCDe886IylqVwwV++iEWOY/yrBS6NQLqScOVjHYc5LTF0CiLq
Eq8AezFzFZJeG6ZxXh4N2LZTvj9xkB3IAKldvFdeo45gDn3RLuCv9XiVvoXi8hjBSVLIztBf7WrS
DB3zueJevbZFa/PzMLRiGjYXurB+utd4bxyA8KSYgZ3AeWMYI4gkK+NWmzi7oAuu8UTK3vELMYbz
IxEcjscpEzxCdCEzQnhyj4aIiUT7C7CFro0a5MrqerZGpOIm9aRgjivB0N6asp/GZ5l+6bBuxMmK
Qi4kVJoqeqhwVXRuZt1lymVMOHSGkIsgb/f83WmvjPZ9VJVadaVCKODuwjyg4fwP4AmA7rGKH4Wj
aQfbqcdJKfB8Hul3nM8m4a0Gf+AJOsagmvAbb2HCkuG6NkUysPxyGZjfXn63clI6SPulex1y9gnj
vD4X/8aal5AALRDUr4rMrGJEAqOV+/DpNV5i+ZxVqukz31RE68BxF5AVnfPBaC0uR9KHJtWnJ3ck
1k2v8ksrs+pARbRJktJFS+9Afe5BcKBSmWXDiYgrXsNRHYpL0DN8TeFZCZjOTecWKhIEp9dwQmB4
MyWBheXYEAd5c8VPPGI5dcd5+s/BLrlOYUlFOCNqrUlfGGqjjVuAImyRKRm++YTfrbJ1gkXKtdG9
Ih6OgTS00D6So+QWVci9R+x17OR1tfCtqOuHZG0doCZdXXVy9kxRd7SYzCUBj1oPJmQUGB+h9DiR
EHspEGxzGIzptjBJzzYYYPlMu0QyId3pZ0uNBSaZPeLEvSmFQQjpQTdEJaF+QVGst5siTZsQGbOh
qsGO0GNKZTwhufKRqtFbzbUEsR4j0hLbdVldy/wd0kXJDgxxdrDF/FFlXIxxUs5Jfqp4+MSv7ooS
MBuU0D7yVunpaETkGLkifQsH8sxhG5lvCQprboXJTIudOIp5Jh96Ym/AdSveW+oqMYXP8tzZzYsg
9zQ9F2MFYN2GV6/2/iCyIgguDapGZQlNdgeMb/nRGccgUYWuadKvVdHGbhKTYKWQOcf3B0F+1uh0
jqmDdvtbj3Fe6wN4563riutei3ry+KiyDSnpXv3WeRwpO4/hi5TLQ+FvVavMlymCrLjqu1QQyAA0
qntuuOaDuOv8fDM/2ubNdF5WhNXvUCvmqaBIWAM2hSvxb1dKkE/TL7/aeXNT3eVSGt01Xe022nCX
ns9CT35V8AU9MNHwI6Hsnep9mW8CnrWQKfH0BsNyRGFr3d+GjHZ2iDHiTJ7yFmt6ojft2E5MocVz
LVKR2fn/i/DtuuRyexo89saFVcw7qKRnSsIUgOG4fpJx+tkAAoSAsGqI4DBJ0CUeW7A+5pDnN5gD
E8+N+crNBKpuHyhRI/w4hfWYE4+N5qmWP35soHEEVU5vfHMWfhPsxwC//Szl+0uOPyG8QvXauqie
zjPqHHMWrkqICKTnxJfuQwmhZnjwuRtBxcoWyVQHqDyDWsAmT94uGiJK2skfs+kZcPNrRznQLeJT
sX+LJ07SDYtDXNK5K9PqFDWk/NbLMIqhCj3G8FeKmzgBjiA+oK/Kc+NVYbAjuYuezgwAHLpVKceM
kz0W4cFqSi8Gk8YVsVcLM0feTZ8PlDMBnweWy1jqg7mrIjPplFaD87D4wJpnLsAfM5Y/45d7l2+8
ruhKhNhRYYyDVgK8zJwd8wh4fD7tfFCjXo3jomaQnc3FEf1WiA1pu80yF7t9AGMpPRd1IodQML8D
yebIgOV8txkld+Qzr+hDXXNBF3kEoxGMUUXDsYQ5o5glZ1VVK6n52hSLwv/7wCO2Bz24k9ihZ6/P
J6SwMaL4ikQiHSq4/FQmsK9Oa2cJtctE6g5AB0hwT04fNCikC9mfZOxI49Jx/PcFd8z7/2dHd0pH
HpYss8+ODr7twjGkmgdy0hukIjcIzF7bKSNcwxpw5wtiCcAW+Kz6iykypWeZsg0A2Kxnr+ZRPqOw
U0+AvAAPS/xbYlK+cdIXMnrOW7eAOkwVzEn0g7L1OeO/hVtMHiSHu1iAmfY+eR4sA+Kxg9pi+E4V
hKOY881Cgg0oC/K8hxK9oyNN+ZNdjjl/UAmVtjhOVwAev3V/7kPkWDCCRG/aVFoCYC9ckBYvVjTm
PsZs8gRU5lbYVPzT3gU2pB6NWdnHTvfoqEoKzTwJ3xhwznJ3K0IPh1LPKQm1zPr+MjJGh3uBJY7F
VYrfAbb4GF3HY3UpIh6g6SrItbLnJOIFHIHQVWHc4lMGGqXWtQ0aqeYLtJurv57+98YBz1MiAl/Z
q3jf2Ns0HvniSZtDRUt/j19P0i66x6yuqaBX8O7BgRChpKHm+6L3JadgRQQyx6ln79caaWFTkd7a
/2H4kengPbVSvg6izVxk6S/BQNMQ0ltOdBn632NXYsNmSESOX0PvyNi9ENr6frIRzWQpesUxVjCi
OXbROlZL5XinGTqlQ7j/6oKv2C4YBQ6NiKkw2n0AkkVu1p1540+jjQV5gL+v72K8Uc3kMm0Lhucl
V7KRWmCdgGyF00VPtOe3sCvaESYVr0p1FwUwTrHZwQvh/6eCCuWLLOfLf1G/AlT5zJVU6DryoWDW
wLk64P1p+ix5n5gxjwcSNzDHWL9PjvAfqNye+tnk163rJOrfuWS8sxB4YdrrT2N9g3X5ayK29M1g
Wyo1CpbrSL+vgkAngo/iN47/QCQogH8Qb2pwIrZG0nsW+1HFEW1h9iHdElduIrFEfxQ8fe6uljiE
tMJscVFe2XK+KhhXqM1yGFJqIappUZIEp68DtdAe7x4c6cPKYg+if+h3XGCyyTjYow9y7GSOIX/Q
1gEvsrCowOta4Bmli8taZR1lVezLqXC19xjXCslKeqRxN6BKxuivDJG8MnX/Zu+Wzl1wyEwfgXfY
Vg+F64ElB4h8DbkCCfU9+Yi0uav9RXAljdn3CDdfRn9aDTkPj1MmPDFt/UAw7Z1R1X3GqdHd82kj
L8/Ifpg3DAS1VfdGJrrbcgT4NZ8dIVp7+YDghyjpWOtu6fKZHQ0H7Lqce6+nsAt8BrC0jvxdIFxm
BGllXYkdLQ2ljmO9ep7ChG0COupWJTyrY/amKYrvbCpuynmweaV9hqy38/KlxhLIVluQC8hSuVC2
nSpzHpLDd3ErTsJ3gEtLYpnTrJxG6kb+a5iYzQLjmI2PLHyWcdbFdYDbgrBTpDPDCSC9hNdJShkl
KIdFRymU49YXfOq7JzQ2VLXmWrmj/YHRMPDSVUMy9p24+iN88p9u7SHs9sOts6btzQMtO2HVyKGC
xVh1ZVhmjyeGrZEOzNWxJ7WkZmQQ4QGXlmRTAYgZ6p63Ug44o/BxdIHA5j3AjO8GVxYWug0UCfvV
UlZGPsM8xBKZMMsu8TyCbJylnUx7k43JwynUV/iXBwMbSCI7N6SrowunKN18yFqYYexVsMtNGt6P
YObEXJC3U1M3f8li7Q2y7EAstLM/Kaj1vMEpN2j2ff5d7T4Fu3MmkM5dBwxr0b69DyjBAWPvjdfz
6LJTrGq7kGKeW+7fVs9ROJLz8Wk9BiL1em11LfE0cV8ZdPuI4TfeKtVpHGHFg7v5+r2kElHhSObC
AnJGYpKDZtlupiV1tFDU/JjDUXU2V+WHh+dwaLCrIpbQbtciqT1iy9No2NsIcqyaPMuMLX8rMP9J
ynNJkF8dDyQNVMCwBkQP+Osr5Z8VNOaNz1uO4ihjaYJvBmr2y54449z5HS1STEtS7YqeKb/AZy2I
Lz25XDlqRo0xLrCB6fEchhZjhgTXgTzojFNQpXU3ugNSM3HRFYTWLzcWKlqprrYgd4GKLiM7iR0C
6iYgUa8GncNsNQiDCEErbmv2/ETdLhl6zzi85cQKFy3O0uWmGfOFA1L2dyCmJjWLmshrTEpNhFwk
mi71zFwy0mzhT5EcXRvEUQyjvFpFhf+cG3Cu9omgCiuazQwbCGmknRwQy9cesCYnzEKNdX9Desc4
9YtHHcN1w4Fzx2CKQciP4O2Cs27xTrGS7lM7zZstOd57qXdWtEC33UNVjrXKgSKs0HOCF0kz75cf
gztEu9rQpWHXZycEy7jP4dhu6KH2mk8Cnv2qh4vmv4FT/9VuaiddCCrj8Zm6s3xLwBrOlTCO7aue
0ePn8af3828GbtloV533CmAM2L5qTHITTudRCzlkEKfaQ3YMrgQPKa6U+5mAlGV50FFo+B+YTfwf
n0PQjdfCGsoOnfJsSKyqUfcewFSRa2vkelMGKnYELXWsD/TNldRNHMxVxCRNOSk/mLareAHZBBgJ
iMc/u1Z1xhofQOj8yehk1UauR74oFt+0aTC6GJBCCWSwU5Ww5JOU1v3bROcWrnxsr94ITjNf2pmP
hUDPsy82bygBtgzew2y6n2wWL8jsFZlgtvXZq52/s9HhAW6pmtXIJ3cI1Zp1WIlnEoYqRdfSnX1k
H48KIlx5ICQeOGHTt3jvotNc90sLSmqQrEnk10yqYoZxpYOUjzAcRz023pX5URTDVQa3SGcSaydy
G/ZstpA1ygF33xS0oPsSDqTNI2Vm7iTuzN9NlV+sSd2uJ75JGEnaxk34iDb4Tdlb8N5euiWnP2ag
itNBXioYu+xFAM+mVQqKI0GrbUPubjn8HLAUXkFirEXIelGnSqqqucsKXK8rBHmor1brdaBNOTeG
uv6fFralmjwuOAi2o0SyB2vVGcbvtgjhfeIsOTxrokTcTqymFnR+aAIySkn0B0BlyE43TF2CIsLk
2C5zLTbISiSeTNlRzQb55nqKxXgVKkIOP3lPv7DLpKqUIZ60Zn9Q+bxC6Mi7WdFKBIqqjTP8ah/2
UPWzohL4/tZmFk+4C1GmUnrQDzKIyZjbh477E79nDsNDS/NJWGKw+HemXIFQQmaWeSxx5FwlvR9s
NggwM2PdBb+4ezwNFvE/v1fBoqwuVjvKx6wYs8uD/e2FFTKTi4iK/PQ2ytPqbqEgubEvTJ/gRdGR
N7v13LTfCFIKxjmJh1kaLazsjni3o/h33NCgFYszG+Y1hAM9po3/q9ySTnNzQo98iQmImBAnIJzS
HSQmF//9TDK/3j45Yoav9mMo9dWyG8FVqyNWeGuxGPjg88VVY/E3BK/jqsMtE8aCSyMK+MibxZpx
lCKqLa6aQ4nIldGVzToyDuPH9koC+64NNslYe+Ce8kuHKpjywxQD9R8+amLTPnaI5uhW67zIZ7V1
hyP+p2T2uthvXjEsookIgLcucK7K0S4ObumJ8nm9vt90qDC3KRkvn8kLPctJEwfKjPprnLpwNvrF
gnjYf3as6sDQSXQYuenaWQtuN5jEwzjD17Wxqq+ng5sL7LnVkTIrqjcEi5cpYNVUsTm9/w2RIedn
dsmSn76RI9P3mqPHvy/8KO6MydGrYS/ZSsZ33uhhTsqeDOBiiaDcxJpi/9K8FIoDYBSQVDApkyDL
zdiugfaP320ENx11jHrrgD67iuFnxF9a4Q9yshRHp1isyeoSnunb2cEq4gfXjBNFdjREB8PzPU/b
2npHFqoPW4/v2cq4+/l5Kh30OslxR0RCcvGN+U/b3ZZz+G4/uHDmWN+3S31f/dDEih/QfI6hWzhZ
t18Kq+GzWhwzJsTm/B4ZFc7Ge/NdnqXt8bSc3Qe2PF4Rrx+pKOrVuIMbUOJZ4+JVRlb78dokkIcz
s5RbL0qtwK5J7lRCu4HNGI211jw0SZMJN1YvFU3V+f4trlRKd+eYc1FCwVTXkz3m0YRXHS0Uz7Xa
HFPq3F8QHcag03f1g5VUMMw/28QN4RA8wboyeVFSb4+zJkYPxH/aHrcVKZoo2m61r9/s6hI6YYqf
p69xkbXrmd6rk45VGia/3dMOjK8Q7ofHhbDD/YyyFinNu8uG7jQbY6ckH4x4C6Yk00zwsDWwsvYT
gRU/gSj1QFrkIAPixvSSkhXVxr30ybnQZy0EMitdcW31QapogCCag9M84ZHoJP22e5r2zfJjKzmB
YFmegF6AW/igvzL2UQf6wP+PsPe19iyibSxIBt1YX5NZQDRUkegU2hDaiInRUGqWFZi63yDHEkBh
6j0ef0OFctHiysUUqQp9xKIdapoShk/wlxPmRM0uBbS/nQp/IlGrmCQQDyiokcEd3GlSED9T+x5/
NlPdagkRr9IXUjLOOijPabWCHDINnOgZJps7/dKyGGDeS7Gni6ios6OMQqt0zwtTtmZkaEtKE8ny
uI8W96CzWiGxUxrQz9Xri4cqqbGDA7+LzwVSN7Y/b5hiaWjL6FMB2E63ogqrXsMMxvVFjGZRn6hr
ZcEa1aWdv/bvQh9kP3D+Do1fDoWoD7UAPkKG7YLWEm0I/9BuBglbUNWcPvSi6AMoI7Fe0WkHoIo+
hzSfMME5Orc5YLtw/9L6IJIONEUUtofmXtatpEjMSNpOWPsNdHa5+vscC+umK6L8/ZlqjT30791b
9bwp5ZYn11uV30hthU5YUr7N9b/TVVIbXHyLyVA+KKLZcnjLmP5TUgkJNBLs0qzkCn3A4lfYOEXx
DtqZcYCI3v9teG+Z4vzFGgnoUTJoo0KRhH39YSka77IUNqlB86hhzhFj4oBO5+wKhsx7weQgYPvA
oT+jmMyyRn/MuxZdXQQ+/+JxMYimegaGOoY4M+diXNiGfRgxH3nRsTbUT5D86JiRnavKCVX6r2cj
CNqjMZPn6UC8myCY5WefcR2VII5no/rwjIh7RaO5LtsCUEwJkwHVUYPmvjSF48IsGHw0JCV3aMAf
6O7Vmuz8Is9WOxmpTBHOFmy8FnHpb2Eycg5w7/5bzjooC9hw0/wfvaiS9ENQ4p27lc3hCSUljevr
0uIf0RQQ6gsIneHUpnbvpJ4F+iEIzmkVjB6fa9MuPbr9xMebjOqTvw144R5v41wlmlTyby/KQzNn
uWNWrROTNMGrcKxM7EucyCYJy9AcT8TioDDZGXpFAi6O0II30pI7V8ggEE0tdXDs4fewfgW0pEAe
/I1WmwWmdrB+C6enJNcFA5qkyXE7qz0VuUi9Jm4kNvJOojOTlKMNtAgECCOVbYNmtYWAaJMhjD89
Ww+N8A2Hzz2qSqu/RNnnC4+V2exSJCKFjMfik927ccafjL+8G10um9MN2dwawTfTgkCmX0HcAELd
CHvjybzJCk4APOBvEJKeflLMz3u+I1QshBYc/QYkgkx1YGNd+UCl7KCPgd1EldrUGoWVYaFBkWQ0
lxfeUvDPNk6JT7kM20BE66GzgYaNT2gb/jFgwiViJpOE3pgAdVG4x34U3zF7j4asKuZWzKailm87
rFyX51XhejCKdfLcdAkoI5PLZm8ZMA3VBPZp+yqIkKIsO7wewg130Y0baAukY0ic1Nxhi/GN9+xv
xB67RAVHYJD4OjyfeNqqYrT5hTjq3lnAke82Un0gHHEYTGQ/b38/VeYrW36cO9eudBX+l+1rMt6G
0MjSa7d4mLEEKmZjgCmTTbJ8VYHGi1w7DJDVbjXtCLX2jQUk6/Ik3qHsrOryAV259QUlJHJtAbrv
FkSlkR7iqBDhMEK0gqhkzlmcXqgl7Dg4cXfod06+NmvgO2HEqBsfi0QpZh8rGbRVw4dqXffS+YLU
4Mt1lGdChmUvht9Q8p60inYBP9shkZW3igHVjTg72fT7THDm7E6y2++b17LOyQpSsjfe4ujt3G5L
Syu/QgjHrqO7VBlYRwSUFV0FdwzvWMcSCdxT0cML8MmDXE0dHmBej1HxNk6V3BQqAmD2D6egYbk6
IQC6DF5wbEXXxbsNaKVZO/J2XjkzeCLtPjwnr4rANi9s0e63F/q5JI8kKsxG9e/MJSERIudz4T+F
cnzbsOFdUonFa65Ow8aPmilpePLndT2WH83MSY/Rbc4r+SJPt0aSBTWKc2q5vqY0kO2/1seZGG6Q
JLWa0J+LPszAu8wMB2CnA92rPr84pTY/fqgxqNdPMMDFfH1+V3eyfwYjKCfMbcG4s4FeHtRuzriA
FsbNZrQh4hyViXb6XSaRPF6hWoLA+57TLA2TUJJeBYgt8ck9MlTl4OtZS6aHF7w6/REks2QOv5nR
E5EHwbZJ+jWCYqATxL+mCiU21AC/JV0HpBzkemqG24WUtQmYx2o4qu4guDCL48jHOjeCRKm9mKSi
Hj82ohna2wIV77e3wqRhIMYZgIvfnL4JIcPpQapDLKGZh806GZQNLbT/WiwYrLLZg/HJ4HfCVt1q
Yp3qZ5OkPGNcerptRHu6hDinhZ2IAcLmSND9+YrijgeBbAQwAKVnV/85lAaywq8ckY/cWWBC/2tu
w0LmycAeSpEhUCpec+rmTFgk3tLHnmpdDdq9ctMMBu3Waybak4WEvfSuszV6FIKgPcqa1ZKqeO99
ApAngLvpxgkkV+h3yre6/bKUk/VvFbtCWT3Q1UxTUrC2yYaWz/1dtYJMjr7/zf6Yq0yYZmjr2cYp
GWJ/RFPjIZQsf5HgP73eBNcIEMmVEs7fdwJfe6VIIasWIgc+7D9Nyp1eenUV7/nFEPovA/ck80EX
cYxKMK6sPE2tChSB3Jl897Ph/5p/QLeKVRuMMs0vWFM7DH0v5flpm1Xc3umyJ2boZGmPgEa/7Cpp
YqzzEz9QbnIyJionblCDEKexMRVy1H2xBXdN6Jrwvut+QI25tyk1HR7GFKfNZRBvhR5LDd7oySge
sBiI5OfsZ5ZZi3C9nx/NPnqpms0IS4Nk+VmjV1ULIhJPhczXURWqbiTwcdr4OPonuiVyz7A/Eq5q
W1n2HLV1GgAj/V7t7mGcrQEn2ZuDaTenDRbN4Tkn0R55wUPnu6J3tGbaY8LmCquP7DWoarziiHZp
Q5o8MNZc1yw5krl7fTmM9w7ydFog3vBHfbY/2cic1/9FB43AUziKH6+r2Wwg4GalrycV83I20w7z
vV7+Mol5f8fQYq43JehGvOvimkZGOedJrcjjtdHiVt4+lVhExwiZ6Ue7+pZ+GRsu2nzTO0uDo/BQ
VBJGr5Gzc5Kab7QnH8TCyl65n8bfaTa+Wa9Z2AiHcB7X+SINeALe7v5tCYTm8hptUVR1Nwz3OFcP
35eYJD3/G5J7LyOj9c47fahdqdnvYB+gaHGqy9K8FZY8JOOFGJ4puD+rQrtsYY4CG/dzcxRuVwKo
0Q+KJNavOMdXEvKswauedzv7eI++VNY7YzT3vjeKSZkz/GsfViuA7ymyjmA3whYx6ZGvaN9h+wY0
XGdE92MFf9esTVBUidl6gSElGXih9HyLI+PxI/lezPCTwHv7GtErOzCh139iZVTfuWxw5pUelezn
Wtv6267R7V72pez7g9/NLqV8GaRYYsCq2oV8q17RpbzAqcZTDJQihewme7FwJEbaUQ5EeLGkKaCq
/GU2/PVe2KZSYP+mWKuCpiIwzJhAPl/925ZaupZgEQXVC5nH4/0StdvyRVZTBpThQ0M60gN+m+FR
QAvl4AZVzw72S/Sw0EVyX8IO2maP/hV9jnsVq7reMm7aAO9OSGchuYbQ23Lh0i8CvlsqArSBIZ8O
+wk4dGnu/u6nPuDbDJ/FtTlHPMIKixDz4wStoE2GRhKYgA9EqgKkugK5Kn+s3hfwuZBHOAenZuWu
Lt6sTjiNSUXpYPxAZ5h4m5Jtec8EuZGvNU5ElmjQXlpCgbbDfJ+TOyzU4GRojguO7hp0HjE6+gzQ
qOPENVsDgjVt0B+LzC44q4sfLpyVG1QUmEaIGLPGS/uPHDT51m02d1oqq+kZS9RtCTFptA6caK6J
qNsUeT/k9FjLAW8mPC2FTTYtD6yWmas7NWDch04k1toOX1YlYikxOE9+JZa5b2Ljt9hHrr66iLy2
v1zyhIPBUtT94GtLJI50JMbGvQBy6ii8yhxv5sTw9M2X+C28f8KdPhwdVFnCW2GfFYppyHQKw7xp
T6nNbG3Lpnkp4iyQPinMXPOz3DPcyhaQ777Y8gKhcf9k52Q4uZ9+tIxWaqwM8odoN1gcBWTsmwDP
yO8s7KlsopVZzgA8LSBZ0pc0aw5Jd/poaVLpC+FJYmlOYlDaO/Ia0wnqZ0kfH+Ug5NxwbsqWTRhW
gGjl+k+EW2WbsvSGjU11apZ4u8J6tR+Tb7RqLixrjfUC9NyFaz32PC0p/yLzbXQ4h3gJGlaAZzMb
r2EToU1l+/0slWuCB+uCnBib9s3iVjtW8U9qnVFz2jNdSMpbI8Y69ibitBIWpvmzZf1rtfqUPqxb
+Ue0r/ZPvIxcTsLOU2bFuRDX0G6FpioO14LrPFUn1Seu8TL4F6sCkzVVFmpnYhv5d86hywUn5rIK
SvlmvFq3vX9dppZvFrrIcHeKqL3nhQAk8XOvUIyskhcX0uC8LCPKfei8tmGJgfZN32KLxEDasKST
XcrQF1DP5aWd509BYlAMvoWTbLctPmd0CqWkJZOGj+7eJnrSP5sz3CxdhL6kemf7avrXkU4RX2c0
NygtZl2CFd9VnB7nz8A8sM2DKMaXhvOi6+UOqgV6Tj2v6AstN+MbThVHSMzwXNxaQ4xDxPfhhMjw
aDwqO88s79joNaHCGLMykIwSuOzfIRW1mZjz2UUdiL9ThzuaKtn3mjzq+ozAX5D16Cu3EdBLU1Mi
IyV/8F9JLuBPccu4Hj/g8E6+2SSEKE9yji5Fqg9bVM4vOpQ2B9gBy/WC5bGuAhuR3OOqx55PVipr
k8rs9C1TDFkt+9LLWeQ6Fnoow4bEiy+qvKB1p0dwtrvj7+viZACJVxXb5in3QFm//QXrw4yCtjKH
1ufWlO5e+ZYr8f/8YQs9TYCh//94iXkaQEYvX6+h6cCvzkpqMD4SwkLpDJlw7Tiu1EJA8cshnuU1
19qtxar2KCkd54pnTmmA5+q4Pb2BaEl+BCEFPm+RXP7dXqSz8Nchjpa+xc6ERHfHCciDeXYV7oeO
HDx2VqYbvdNMjhiCQ//fiyAzim/wozw+gRdQcWTwKKlBRi03v//YCeJWxzo9dlQ8ibOFekm8hGkE
U3FRG900wSyR2RaRzOB2nMGjBb/rX2Vv+MOCU+QF+D3AhWHh20mhtlMeP3r1p1GOBwY1tM3yAuEE
ivbEgmkLMhRCwZEsQdBc2uM/Bu7IHUhftLM/0GX9oq/xpy/ucT2JDIxihki0581REsm3CuK0JWGR
VgJgB3U/0P7s5QCjheHiWINLcGaaM3CMrVOQ8+VSO9emzLej3piDa6z57/a8bsYD3+ov91MwFWtP
Xg7cUSeA5D8iBBlXhIQz2bQ9HAJy3RmN9CFcXTZYWR6YOyYkRlAkVymdfzlWhmIsCIIvRicdWsEK
lwl1fJC2bvCxVU10Ia4ZmTws9srrIwC0/lcdYyMxpVK6UEg6qrVL1/FNw/saO5H+4DZuYK00jihJ
xkH4S8O9ix50PqCrCy6D8aXkx1VphdDFtRv9Mw0A5Zu8STqIzY4Be33XjrtC8pM9WBrW+3mKjHIh
ucBONsvDWFs/Cxck7Zq36XfCPbi81Cy7mL7bv7lJ1P7os5NtHv08LDywb6yNMQrIttIKWaPm2pR1
+hNLsQP7ZlIG/65mkLgTais6PEda+y5oQn6XvEIrKr1Tmp1vH+Wu1SLNKe+fOLvg0x8MhJCqJ/l6
ToyRJEbm64wOiYDg7dnpKX8PQ1o4dAv1LfCpOe6MJ2iZdvCbXDqdD7Xzz8Fdtwn2rqGV44+2gk2b
HcniszAETCbDD3aN5Fy06p2JbQv3d2KcHvpLvjlrP3QwaJcHGdHPvLa+1SWYKD/cPJRMX7wI5vz3
BAmlRkS3MslpZO6bZLLekQMdf35gHak6vo5g+zI3gAK/P7Nhye8B2QoqfgpwYyLF/mYqyFGV/euV
MtBwDtbhf2gXOwErFXMtyBijRJwr9csxibKY9uzvkeTh3iugKMtws/U3ocwRIZ94FZZQGScp4HDj
vvvIRTLEodeGU0jtspz6VaoxrR0PSbPRy185dSCYgB7YKovZLolrKhnNObY0E9ybc+zIdo8tT1J3
GW/Eg51BxDet1phgBNXz1VeF32fzCAMRIfQjPFRgYxZtx0q+8Vqoog20A3Bm+q8tdy+Gu8i2nHjL
ubfJ9gKwEIWdK8V+fHJQvSsMFptUzyzWwZFNPCfk8CLvdpdgkfa7p07sw5+54A5sEwONBe/L+mG5
SRSpjvLGuNrJQ2P13q2NRZqPNK0sOzvHhsza6LyLV7cb1ef06RF0TtGXej3SxSZLDFttwi6a0jql
LUYDyZQ0O+TvahVECZLwi2zewETMC+gdVbrBw1RK6n3cDf2R/9Cyp7Z2yRkpwJ0M9Z3rM2rrMCG9
Ro9jBpWmXCiqgaAYJEytvAhkr50QpqtCDUV49Nth12gdvHF7G9YdnZGsibEIPS7XAsWBpvT2jrH3
q8IgDmhXXPpD86fb4BFOsYn/J59SYQYQORJj5Y6FzKUmG8gsDKNYvfYNO+3FjoScON+9muAIy93e
9IqBnpmtx7APsW7YNMkFEuSPlr6/CXoW0nebidp4jda3d9rJum164deiAxxtmgNEzoLqEAVBzdO+
miXf+40qaOWsX3N7j4UtEiH7Fu4Q1Q6hTalEZdtKZbre7U89kQq8SewGKYdUJBNEBBmf6W1L48pD
R9sbbt2qcTl7CnZzXo4lcInFhKV4/eZ0rA/3tW4OTMeT04emkhOEMQyxjD32BP+J6m+fmt7mMe9x
c5GZ2b6SkshR2f4cbR53YccddZ0j8VLUBCNc+5lHePAI6qWDtHIO5rrqHBpT2iodu28DEHUaw06W
79a0sf7CR5L4EW4ezC9MY0yHVz8HpnIUbIqeAagcMFqtUML0FgMwfNhcdNiVHXUxkuyOZRb0CBTn
GkZ6mqequkew0gx80sQUIjxeBhcB30jod8isV9rl89HNeQmmBR3k3An5zLnGkPwOG2UnJ/oWBxuG
EAPecERmvbboenSrbactbdwGnZIl2C4pYqiMbq9qa5IAMunMzFAfPL9QUlo9qOlb1CccQGzwoBV5
chgj8iKm3t5cWJr5Qj0zlFw+tc0MFxfPCeJv4k4Cr2SJ44I0h9c+97NwN0wc1VK0+oyrWjYPcsQZ
pwMKXKwzgIwrNDrFrlK0qpI8yvjcJfYyxvsDlNmWfnQa4X/drtQBjQCKKE1Ti336NICFDmBQwImH
DNckl0gsrTOZkM1fxVLOduAAwBVer0itPIVT4L6KSuY0WCfLung1+lcJiGtnGb7WrPwkrr8q/qR5
MEzf3YwoUrVX7fB91FM9CZ/WKivs4kix5eO4obII338N1tvZK0Zh3ua3NzfcTtrhqQEpWQ24QJEH
MBJtDqBp6jHX1/sMgQqdpvy9UBgZE7mIl5PtsUND2e6mlAWP63UNQ4AvsZJvFtvyfG8mLdHze6au
SVleJWtC1GIc+JqQQVuMnfamGTyKNz8zksz5v/J2ey2xQTCoM3g8Zx8sQboIGnvocelpwZVsjBeq
yNqdSQNjqX+StmMZz76GjX02AedPLZ9QnkS5HL5niHoDJ1TfJPLpUrJSnfjTKKKEOASgc3wVyS9r
ZnwduX3fS6Kgfw+bOrQB6wW/D5lJOdM/Wdf0zMZPCwjpvQpVZu03JlCgwEdeU4L5TRHo+hMe+E04
tutlBVMbCohYgH2HN6L7A7cLPyVU8Nh8NFZ9PxWiNstnwOPuLh+3xKAd6x4AqzMT3QlJr8GxqpJE
V65FIbUoU/LzxCu/cxmx3FIUZMGhpIm+ORcqFfxEOZMC07tkdPBAoF9IO6rzFpe/HP3oO5hb80Tt
wb7qYwNI8EjrCFA55wYG15cmD6sQwSteb2XlhV+0aqDq8j66r9VWUw/WrYNwHuM8c2W+lkFr1MEV
YCeyAquAWWmnWvW4NKM6ixrUIF07WDmDKhIJWhxgdX0+RBexZ1DyJupyNDQr8Da/aYpUcLEQMeG+
pjQXULDl7iWayCzccYGNQ+ldOqLRpZy+/aaZwiSVzkjGyxRVS4DjeoEOHg//v5PY6L0R20+CmN2V
WLAD8klCTAASf4XF5Oa4OJhZeAc42eu9gkbHQKD2ndAiaQ4W6M715OEvlREEeOq6yfUQ3vELRw2K
3uWABd2VzbbL1IYL+osH+HAK+uouFIRFXMBl3yHVLmPHs6bcHUgcv2seIaldXISCwOOpBi4L2Nu2
6CuNhJGfDRf9or98WgR06p2Hk87AV3HTk78tuCDXCTK/KBFYz2vVp6G7ck6kdR+AUcT/5QoP+1XK
2ZQMDjyZfhuwamZ/eZoAlkUgzYQ+X9rvPu/nojZtgM2F9ufiXEzH2dmZj3epsgKJsRl7Mi1Ao/a9
NLJdLhA6zd0/Qo3iNoV4YldiEWUzpFoD6sfm227Rt985T9mkSWDo0wh9zteXDde6cXly9I1E6eIs
qsAXarGGsYbl5WZ5bVQ9N8aATlZOW/nXUUTW3pOGqJ5kHPJizUwZnEKQK5mTgs6ML4Upbh6q+vua
mNwEgy+VGAOsAskOWGwAG+48+iremA+A2j5yzo1Wk6zoFK3gkkgxUchweltijnmWY3GCUNu8uom0
Qo6kPN6LV8V/krAIRfYpcGSPFnWIshZp1EC3C0N4E20Ix2hwZ8rNE1LnbTtY2CAdeiu3KLrKjrQl
kLCOs19psbGZISzOZHgTlKYalfYlTaLvw7+HFK5o4U65tzeDr1YOWA4RoedWmP/lRWmsI3mVFr2c
nLJll/tE21JIziXoRdhaPm1hY+t2V4u8s7i4MWR4ew4/hKYwDYOhG45ypDxn/DVCYel4e2QST3NO
oi8RXkQbNiM5lSVoExO1zhj7ibsvp6VRiW++Oc50kJPdPmqmO4tYXtNV3vfN+bcea2vmhPhF7vL8
iwkSEbXANnHX+wvI+McXRTlzU+eD5b2qJ12HBfuoKHX+txeg40eYN/6USDQx4jh1+Q7Pg5C2AYnn
Ot2lwg1N9N4VNRzBbHWmdrbZJIPVqdTSE/GB9IiaqEKlR0ACtfBgd4DNk53nPvboKzfs2oZcrx4R
ROhcZWZTyXYNkwZN/xvfZ3K9vRecytVApZmgjDtIMV8YsLWGiuhiE9w8faNw0TyIlGkZhha/l/+M
WMvqlFVVxSPyuAHIhGLo76Tlk4PSW2k0ImK5L8hhjaT2y2oyRzWkQ5Vxqym7u1yYfDCepIOlsTJP
MQk478JmbexmpIJHSEdfGv4QXDyD0xetzb8V5Z2gz5L1G23AnuHrQAcEUUnBbw3CxqBEC8ouWciN
y5bVzYDPv23uSlJ27HLvUmPDIWulxvpLzOSYah5B/HGByNmcDqHjzmfbSLWcsdFqPG3UZUzFO9y0
QYD/Yvmv0oBoxV1v+wv6Pn3O1824auWPOkWxLlSLwVAbbK5x+R2ghOIKa+RBCtVikxzei3pwt6wa
NPFtpYE18zvL0LKfFouYzxqe1NzUa40PHjRES+wbJp/Nv0qJidJ7/1ZAYHmnoXrNGE1uc1PI8u4a
rTgp3NdvDZX/TtCOBoBffQuSVNvTw5InjdNAS40nw9vn3LMM0E/cSLj8gPOGoUF/ZpYPOcx8MTps
4nsjsH5uuUOyxzYgulTtT4qVlyA2p1GLBNDvVqkMBAW4kMCf/WAlLcbQju55LqdxIAh6hXcKMA5W
RC1HtYdYYWzrcJXWh6QRbutu/tqSkjaBiOpAsN2cnzPUvCSXyhrJfqtuc9mbocWo/XWVBgfLjCAA
zsByQhGSayFhu3iGdlstAFbu2eQPTfsw0xixMYCEyRZD/bF1FPKTGI5iYw/ZXltdGyCdk7sgwTuA
+bVy+SriNLKFlG0JYIp5xsSyS1fGIXWw0uoHWnjbq3ldr93pRwev/b+yGe+prlNZmXsIeqBwyX/d
XDnTeJ0HomKLhG2wMiBFhe1DEJdOIt1nT35usC+jEVxTagVlOw+DC2a8TwfqTEfYkSnwCA0tj/ne
FRchr0+7Ozla5ngUILYSUwR15AFhBEhmBRHL1Lts1Pi9wmSy9P/yLly3spYx5yhi4GgBVGVYsYD7
BioXMHKnDdBT3ZWTWad8n3pUhEAN8leS3jkTGJDlTmfX/nubBQ1J6dHjDxQ3VLangR+sJzNjVSqP
vJQMhoorWhdsVeoR0HWq/gmn6F1+FYVRqXtugz4zAvlzfDCRJz+jt6UM1+r16vFioJww6njp/VPb
GqskS+MifVyXZkrtMjhfQjQ3lDNkfdaPc5tW4Akvxd47KhxNS9B1MWvdxQ3O/nk39HRr7f3TWmYz
t15bRz2BPLhldX+9zjr9ItkylCYA9YC5KfcHc1mcK4fB6RfaN5iTz8JzGvK9jh37Pe80Z38ynxJ1
dOmR+0qu2OsjsqNDt4Ga3YGjT7rwufG/QiEOCrH9HCclg+t82pWkYgcF9ZvUXco8sHHQbR+YIZIF
rOVzT0u7ZbW/J18fadeKj0z/u8w+HhXgzgXc8MHqFpNki1mjncJymFwtNTPkDGWbKXtiknrQTMTa
dOXE9MqDRAhGoheW9O+yJXnm1Gr+3cAvB2E8EIToVu5g1t1BZXkcmMDV0Shb4/f8AlN8OObrL+EM
kPPldNlPJnj/iATJ6UHMiomVfLPp8yoadCVEJ5bpDNVDEtlrkycDW8yHDLhPBwpU7ScR3FOro7UN
sTEb5Y0I2qtR/3YC0QW7+J7GqFvhoJgorCDxhlSa0z2ZU1yQkY5XQzX3EqlQksewW6h872LORV7G
yaDEYmeXWtIc9cC4/88Q6X1cpu2FrsufMdCg5dBZESa3srfNmIFE6tfh42eufeMNrE9iLojinboC
PTho7KvyAs6RMfdh+q9hNXREATVvkDb3mR25B0SrARjomvJrezgdcrVwnL7BBBPmJ1NoNHx4vrDb
/2zY7y3BJJ3NPn9Eb8+EGLyvpAhlG7qW/xzC/SU/PPwnvFc0KWWJV1v1nSTnP2Vja2ZWVnPJJi7Y
foaM8e0okc/gxDIbUZbMYwY3H7uVJEime2uvleW6gguVv6WhHCww+L30tsaWQjoVjMYddD32QqA0
7eEdU4p4TxKiusBjepSSUiyETCeGAUo5POPG7MjYP4AetEcAqz0otdyv2koUwoUAJUffQRJWUqYe
RqVxzsvKw/zkUOVSJ8vTD6RQWGU/2npTnl4bhY3/5l0LrjBXtQ4uU6Lrq0CF269BPi7rs9TzuTSi
6qKAKbE61fdspf5n/yiX2eVG8lEhGiULRI9Z8ejgae2CVwpd6WKE2zV0hXdinJ5nuxkqMNLjPNnn
SYMV+uYG8dbqR4RQQfTIvVhnBEjIjb5Z5uWRt7wMngMRDgkyB7aE28UMe/vZSjhtKYLc6om0vz5p
3X5Qp2D/gqkhqH201sWjppyKuLKOPrW4KOHZM6ANH3MWLlQkXisxJ5+Tx5hlx+gdLGrad3WSCm8f
ZlS6Cli17PtKapr3AkSFPXmXf1A4QBI208nbslKO2/uTfp/zT9HwD1LSBn3TciJqxa201TjVOwkt
V0flC/4kTvHfrjBjO1IsGHjU2fqm3WGIhTY2v1UJREujaSV9PR0T7NUmso0YiPauQzRiTvt5rypp
pILdh2FEM+TtQzveU1j/B5xwPiuJezuJ8W+pPIzotTwXY1en6KlSLboZN5A7EHePQxW0Oq4hrvmC
OUHVneuxMGLhUJnwuyoYE01mfLDU2XnwkySmjh575C1dcqbFg0Y//WK4WR6EDnihr3u9FD9OdpIN
9jJk0endNjBIQSSoc+3RdnA/UWa1EtKAQ51muLX9xIMWWhftsI5oxerg7zLigdWLRnOXLR2sS2Xn
lRstSW7V3/3NUVSK1HP7UJk5pGgBpGtct/YPVD+y6O9hZQ2zlaqA9+Q6z0Fxc0oK0eZKmZVKKBQv
wK+B0iU5CRZJw56d/6CZhNHchn7lhzdpHMHjwngulIsLrWPEa52yw0FG6674+yFA2kfabOpsTV0o
VC++s95mccfNWMKCa/XThXgj6LRQ3oiddsryBxrAGmTL4V0QNej/AbhPFdGaOHmRNeA45lvdPzCh
UkKxyDnWioU09gaBBy2jYRQhfYD/41EYAnm3v7sQrKaALj0p3tPsP/L4qsu9HVzE1Mgmx5DTOaRq
TeJM0bAYkaTdpcxKb7yt78G7BMAwFLXytC4tSKuIxebr2NwbyZJ0lH1/k4MS5OnrqGhCssNYuBhn
cZ3pz/1wWgNSMzOmDVuNu+rGK5esyOSLaP2jidDwW+BPHAa3xXQFrI7oM/KSEy9/emrKKk1rqi7Z
b39LykKq1/rmFmAhKl2MYXAPN3G/JLxVegxu0lzApuaH/giKI2nmZAwXYbdEI8rfXzSEz+mov44w
VJ44dJ5lcboPPqaDeJOz1x552PpZvN1qm3xvOjxadXxXc3RfjWaXSwURyPMFd8MtlSZNlcQTQky8
OAXOj26VHtYW1G94n/SFmPEleVpNkpCDgnN9C+SB2jHWfF06V3JJvDmy84xbBhaVA4g3lGisaTP8
R2VyIDFV0Gkcy5wBMa7I+DHMFjT/ZFdZk9xpIJYcYR6wwlbA6mlXxedS2pwkfV2fdwHHU1oCPlUE
lxx7IdslNe2ouwBZYW0RDNtpTfuyow950nUO5Shq0h8weCoiwbuxf0Pl+hfzdFZWI0Zdv4H17peV
shYB/4TqOjnTl/Yuw6S9+o4pAqRduXsjVP9DdyJYX/DI9iTU3cxPbyXr15jxLHi/108wRHFRejKC
dALwKb44fo05O3tE0bDIENQ/BRMjl/EAkkfgTUobzYsBsT7QQwqd1Buj/5MG/4aILrjeIbMmGNIh
CdSMlytCxwE2TL5Eep3V7h0J6fi8j60LPhNZ7r2lDrB5W5AB1e07q0pweij9iWDNchwVKsG40CVY
7Qm3wuO0DKLZvrkRcSr+byKKUFVLbP3lE31awHR7HTFO305egELWW2yhQLN1UDBvHnentB/rvZLR
eYEQtWlv3Ekor6M6vBVYHqpmdbHs46PSXKz6oRo8plq0GvjxLXgwCRZYtk5eLqlFz5AnJtub1eg0
xvqEBXSS3or6j8mybu65AWir2jpTuIS6AKZPMZzvhNgxzejSMn+tmebNpC0tD7Gv8R2PeguVqUMr
euPFXlubwLC/6bIlA2OS95hLjwwXIyzyg2EN3SCtHKehYc6rpu/foBuJI6HiztxoF4gSMO7EXqvd
YW0gbLF8vncVss83tIW/9v1hcxHbS9MtutB1gC/qBUtt273FAIe84YuPbA7Pg4STb6+3w56+f3JB
PaOp9twjZXdt5Xfr+uiwsUoGyV3YGXc1rgnowDHj/u3tTytrav08SDYBp76XY7Y8iR/6Qiu6hwyf
hyhQK2iCpoCgzurqs0UnqeVmHhMfs0lueNh+eiqAM/lSQ/6egtDAjy/vqGGeHLHWxtlumZkh/qr+
NwTS10r7TzDef/Al8QNHX4bDZl/j66CRGkqy64mSk6BzMCfons5fJnAldUcb2cW6vNRn6PgivcCM
sOSWz1G+d9z8caIDZdatGp7ZyiyPcF32PINhBUjdB/HhVKk8+mcB/R6QxeGnrGLZ1VMkWMKIwR/+
ZVv9SLFciyWBndXCK66EErFswanUrK+YxmUi5nhX4KK7sMnPWQfeZ9OCY9edytkcsVXwRauUPT87
qa2cJaS6XRHR1JESOwG8gtv/IU64vvkxMacGpATWzijVk7VuzXx5fzRZf8j8hTO5b3V3bA+29JLu
k8aCpCkyhx38qLeYaYCw/Dn/sBeEx+ZKWyPj8R4RFfrVYtF+4KiEXDuW1KWXu+EGJ4mStLzAJepu
D+tt/UQYFDg3CVPjDsUdiBK2Lyt2aXlr8iWLMFfx7fuJgGWrNbKEBm/vXWwm7eziW3sLMeuTSgf2
6yiNBIGBjYHQPKBQAdQj6NJmSfDq2s/d+lKbWYB2M3WWi6O0iwz+BHhiB65b5JBm07CW1G3NyCgu
ytiKuj6Wu15CeygKMcrrmMl7Rs+woJ4GFJKVdSoGKOL39bBOxutt80HFeOPaNDrO5Oj2qT/oURGk
zjKWVr7VLfmu/bHoI7PIozvFCwan5WQha5lCs7uRQhP54cff57A97XMX8SlGNFTXuezwsDqMICCv
KwvrUVtWeAZWtXNOruQkGuqFoeb/mYpaWeJJarB9lz9ZV+pWQxATp27bvoGLxxOsZBeiUlyasJjZ
aLX+8PRoByPZjUDLOR//P+CXv6WSpd5ig/9OSHfMPkbnrAZlMgdrvHfFxL0dE4a/KbYyxPS6TsNM
h3D7cgazOXDelBhYN7P3azDNxBFWaK/x0Q/yk1uUNtq6P8cRYwUyvPbDl3R7/UTivBFDaOXVM0CP
23QlInQrIlz5Bf+VBX5GuNdkhhc+AQSwUJxPH7RE/fKW1Sdg7p4wOKt8FQqVIQfn2e7A54W4KI1a
uV469Ra2/pfQ+TZqrOKBe0YGUbtwUw5LqsO8/mGpIG9/tIGNzqiRbGNA2dXE2bnneyKS0cT8YbbX
CGcryDRZXlZp4nxDxtOIgc1IYAULD1zR5MM0sIxeCEkElQJ2537yhstNhAdY5MfmVbDyeZJ7tlXa
jevumBCOndBLaaEIjwoaJOK/3AF5uuPpiatrsGXPflnw8RJFhewRqpQPW1ndTzPwvI5LgZsYgAuY
nUTzbhdRm8GeKiW8pwXjmxznlyupotnSykElMreq+Mk2Q5eS2gJNW+4r4CzeWG3bivZ42LjU5faZ
aQxWRzeh2p3Zh+nDudFzLOSY8/zyvHQJ4AYBx8TYvBbhi079nYrw6CATJk0TIhoCDhjlP/iX8kng
hX1n3BSkW/CgxYMhytzVM9v0GCtm5quAglJe1rJ8hz4Tk5IAVfx9A9AroxlKW96xr8gdrmYbv2Yq
a1FaJgXPFH4J3kwP8VKvX8hgqL7t1gwura2Ax8n6HIJ+bRnYEeqh+gA4/laBdwlg6qxdFHSYHf8D
2MfJEklchQJhlTLCtPxBhoGCjfd3OHtXn05JqwaTNkn7J2OJSVuq0LAeW49FS3ss8obN4tHJctTG
JJt1nUjYmAWeFEetpk5c4ho/zUrA0C8mMWgF7A/36hxZpCi7urqbSJ2Filc/exW7cgFUaQRj6LKu
EWaCOqXJwrZhXnjAc4MZV736PJQAsxcq2iyJUQF3WSJW4fUXaKiC7O/e/NSdjygSIWeqBkAhkOOb
p12JJMl5Dd8SSVT9+DJQWorlst3bsrmHhDB+LvshsSO2CW5HBIcaKBC9B0IJcY4NP3ArhQfhbLY4
6KSG2EMll0W4+54dBihy6nch8l2aj+/6TQG/Trz5M0oWeOf/GkCUvm9tQZvbaBH1sIlrJ/WjcVpG
ODxrMxXW47iS+5UmH4i+g3Ud7oJNt5Sr+0P+XGioBa+twD9tgv739WDS6/s2ZzfGD0FJxqTKw1La
af3oATL+PqDzF/tS8qBcVoSdlkHToj0X9v5byPoIWhvlpPIfI6yyJr7yQhduWSAtuzHYuezlRav1
tUS0MBSGhpHEIB6gzqQVfgS3Hlri4FP/ELk0mrWx4wbcdSvgJVT8Sa7+Cho5YQgOZmtIRVcPmbcq
C7mnK2obrkMc/fB3MPvroZV+Vn+wYTdoI4tNFD+ZYVDpIEEe1Env4RrquqIt5xbxmM/J9Vkc7eBD
zM++CTMLmGsFHfsXOOk9wZZ+EmhbZJ1FWqu4nXLJKl6qCZ1iFHdQ96dwjf8dPj+H9GDnMnD7IDc3
X8Kv18hVliwR7tq84XdpJrXMpr5Yjf5AZcJyjPGDPsDMx4h2HRivBcOemEnsT7fhnSj/rYioo4QG
y108j0LKGujLUBbvznSCPNJg7q2HnG1C/P80GwkQLNvg86WpBmODT+/XSyv7CFk7YQ3hA3qOq6yf
W1z0P1h5bwzPemA6nlwWzzhrfD7DqVXDyIzRC/jAB9uOzdacFfh2li7y0p2gyDp5X1RSTcM4wt7Y
yWe/3lTXmF36xRCXigQfk9meWsHLCe1Njgj387YXPZjPUcob/uMx01JTSoBk2b6MiQ+8i5B3q95I
aeE/NN1NW12CvwENyPQgXY4KiXgI03RXjuWA2tLJaTxMUehOdmAAIBQC5oXRpZbDWWByat6cWbGb
1SDxizL/IJPRR4gyKTgZWizj8RM/bieXXN0KRLu2uQ+4Qr1PzN5E3urUDojBk11gtEGTgYvayeyW
x8plb07F+0w49h1d/2HPUPmccP1vLu5Jl+k1tmTpk5Tk8De9o7cCpf8Afxn2CDeZ5rcYi8FZYo+3
9EaihUTX00axJmJKVmDGlK74V4PsvfMq7/+8GGId2plblGkX6QfxD21YnB9gXDAR2NdcvOXipNuh
qq530zu1XzZdoJmannLJzBg41vPDh8M+GPyeUpL6lG+iDrrYdYr83ypxnaqkSdoTM3GeNnsvOhsk
Vu7/igsazEREK6YlKUYVdu2EfQ0MwNiNCyTdKUqDJfe5qlbds+PJ6sbnoTmstMTNpiB8UWiT8LiY
4aZMg94W8I/TOT6t465eBaAMVAodge8efRTgjjh/ahaBeV/LjcGe8YVvW/ySsMyWrJHAXJUlea3D
DMfyQJiqCgHMpyPWdh/Ud/+9jHNlfzY81Q8Ax0k6EYPuNSrUo2uZCCEpLCb9s8dfYRxi7ozAPfF6
pvaiAhGGlWYyHc20wySXdfMilh0lyWIX3R/oqITbtXduBsR/r+nUuQveQakzZTkNpw0i/F+cXYW9
WkvVyGUVbxFvAeQCCjLdoy/tIZ9BJ4zhucE2xHHGSEm7I5F9hFlHf8J+DHkDyitQBpgqtTr2+Y4s
BcLz9VO2YHIPQXbCz9J1vNovUwGQDC4AE/UQLmLgVdAiqqDGD9b2PVkco0lXFoFG4QZMBDcAUqXn
RYBzdcytamruhj5IFHKlzz9yX4gHEq2+zpIbW9/cL5+bMOXVwb24isbQMYTYsdXY1YStgkX9kbzF
qIwCeWdt8FvS0+aEQ6NJXZUkb9V5+j4NSPx8eBBDbDkKeOdENVNr2fO/pWkanKSpdQKmFyDQTYWS
DazHY64lwjFKKaTTJFJ29a17ho2iMoaQKPlO76uBo93BrxjSqOpsQKg3Ho1xF2niBhSPUTqf7AW3
r1zJbFkovY3OrgYl4Z7Kstcy7mgkiL08wPVCLG/OGXGCdWQP0baVZg919j3VQIEcLjnBPnATHFVJ
vKb2PtuljUw/qFdScB943UlUrmVdGIVJtKimlhpyfZvEgQqGqGA8ZKE+j6bejoimphKoalU7zTin
mVoT3E047TzxJDUDnA2i6kO024QQRKSeuidMirlxJdj9WSeCqyUUKOOYRBXFC8iTrEIvHm6kmxuw
O46oTkd2A1oQrLNKsona7APjadNszHX2avBh5sSfMD6ghusE9qB/6DyK6gFyqQMxxLcP1hf0yfCA
fAM21eASN02sVJYpvME0QOVelix9gz9zEAQWq9gLAEtgPEhzBudU7StMtq0o58DOHeBM8loa80oH
X1AkziydMSwaF7KgoarkUiS+YmH4C22u6Is+jTHt6Ar4fZgFBK0rYE3GiQEO79HptlMx3JBYlJjw
TdWjbkmyrNwdRiQSWRUMwH5WCS/kE6Y/7U0xmPcOgHUWR7oMs8PUpDZcNDeM7WZHGAxRkc/TGKBL
XBFA+V9qOrj+J0AxcodSC71ku65KdwbhXYRShjGtWsH2TKfYoBsm2OuL7Fue8piWgOvWuS50nfHA
wTn91+WAQj2imcs+ica1PeFsKuPDgtsCHPu+sHi/dOzVR+Fditge1Lp5O1+h4VV/vRLU9KtQG5mT
0ehkDfPGobVTW91i41gQiqQI7HxMFkT2UlM0ZBHk7KMJGhduhNDu0ih7WixOr2hknAahtzZXD/7Q
luRLLxyZAthVPH/rEws+O0yKxXyB0TyoZAYdoZEuIUNhhwhP86PoAmdG2xGT9jnuVH1wB8QAqBxL
Y/Cyxuarx7X588RSkwixyEWOlax1bKix2czIauOptUhjvix3NuqL1P2ncyP0UgIc7ZWueIp6qPXS
QHzBhyR28ZYtditSed23a7v3eO0BcmaZSHRTFZtdQuNa9tN/Si3FKGhcCjPIBseKGZjuo77JoQ8P
rPoUy11CoPizB8CUG34c43Phu/lCWbaH/2cFWdZwES6Mtho4YVYl3uwnJhTDFd9Lwr5TuN9z4eow
EZ7YMpNZNLKsApsE/intY414hiMMvZ/gLNFR0xOphVyxeYABh5m1CltZJfDB+er4ksXb+LpSvlHb
rpv4Lpq02xo96xNQSs+U4dXAHQ9dIsyj9Hjl3X3VD440Toofb+/gAqCN1Ku283Zk1koNZwqVD5ta
zEIX/NjBswTBBqtMgxkAaaH4fU4KB7/vzDR7SXcEO9SSoBz+N/G73pbC+wqMg9HaE8UcBZ2q71+W
ya87YutWy+YRDCyOyywa5Lh3+frKz2NTfMiLeHSKMWWg+gzC2TCSC6eSqTpwZvA/DcnQjy4JeqDM
WvFDT1Uz8vY2s1G2vjQH26wvDi7+VEmtarXPCKUVRvQsZcH7XGynjHPUYDdZLZdolepA0hNZIGTc
dCT8b+Y07+KdK4FPq5sJoSj/iGiEY4AkuRxU+8SYygD/bzx4CTxMhgDHtFWO2GZx++1eWxQLzgrr
pqXItB2CVKCUpiPkJNdQQXTeISQlMWmnfwHruP8DGi2TbRnS8QwLc3ljfsTiTC8JZFxAcVUbPqUq
sg8q/qqQBnlakqDzHx24G8qulnmt2+1/ia2JdFKYg7vtyn3hjefgIjLaUJp9CvPaLkHyIrQjAR4M
fOQe3ZMNzTXWyWswYnqz2vnxPLiDg6UrkZ8ZjivLmsvr36/Ev58ZWfs2FPoAhFTqM1+nhoidV9T+
nIb8C/7zOdPVfLLJhSpHcMXd7CX/2g0Vm3muAQ6zBdyL8jfWt2Q7wH0HdJwRAC72rPIsz7JFLBwm
vEpRvCXYn6B2qiulCGQbCIxdGu6hNeToj+nAl5OVqpCAyCJBik1XKFluTCc8W4W3zAb+EFguBt/x
Y26SNw/sUVRUl2qB8A8mLVhzPzRrChJ1e/8pdglklQ40b+rwqBovI0EQamveYeFMgn1xwLx9K/A7
mbgHkVAnPQZIXgMRo6xr3ILmXjKToPjF6bxx6sWQ00xhGM7oQ22AGIvMOPIKz8IdvpHzKNr+DDj9
1/CjvvJu0VXnNlrPp0qZjH6nc4Zh2KjhoxK61TytwyTf9FXc28lXly9EIwZ7kC/9T+jFG68Tp2ij
oVRyeRiPrk2oWdi8aGxn2LwIRjIymam/h7yfK0XOkSp916grUcdi7ohaDKl36Pi9UscMl0VxAmi0
RkEs4aZcCtb1b5rlFwVIlSzFrZJtW56qB1EhS7QLrdzSSOnxpugChSwAX7HIqHbZwRF/oxOc25Ri
IIclLmfGzuQCtDDzgY9EeY+3MWD1h9vNKhJrgVNqQ/3Gopoc5H8FNuvVcssmPqxC951bKYDXrwT9
gtpjdkBJpQzHI8JQDj6zxbgFVGBBZSWq1/dMnOx368Vwm6CO5BiLONvs1/gofoO5G1aZDhmEpOY+
EVZ+eCCT+dKHYjCaIRmkD17SbM5FMmDLYU7+WzrXcgNAAQfHyhe5nYDzGUB6COKPNOO8N4ojnk1V
4urmm1U4XyJHrRDP1X1mSCapeyTkspumz+9kcXIPX8te7K+ELHNeZo4npyBiliSa7vGwdwZ3gfVW
cswgZvvH43Uz956FsYpXjzNsT5Um+FAZiV2bV15uyXpUjmHwFIqzlxekMO/s3w21vH25dYM5tWms
+EyGDM0h48TIOD/+QQraDx48PkQWalWHBMqTBHFNn/hsjZoxT+hX6iLV/NK5vF6/mRqTElBdLqcy
Wi4AVlMC9jKvWoeEWEqWeFtUXqWmXDYoX/afl+6+8eR3VsnwtQhviWYeoSGrWbB7QwmmYvI8j9YU
1VP/ruvDHZV8WLv4KeSjb4zdiTF53Nn2ohNLy6kLJBYcZB2WZk1eTiWgDnllepsDYIZJWEEnwfA2
wEn4CigV4EPGFA7UO5aR7POOlyE47dn3akgNc/wL+dvCvtE6sGLi9PV/4BNCJFF/EUTunbwqUlDB
rXliYhKo91nUDXkQnvPTExtLZZ+Ge+X5MHRHP8WCaiYVZWaSwz0NLYwR8E/KvdRWPGQqTET7Ii2a
a9BvTku6zm4wXz1JKbS5/q5wAyS/d1d4wGK6EopqnQDqtOGtNrTCaEygYRd8DCFZ2noF0Cro8SC4
8q22s5ZBHhQMVidL9M4VKJe9aOnEjXV76e7AaGXQQxM4+vhvzDNZhDzn1korhMhguzFdkZysKMsW
US6FFm6bjdV/bxisbEauZtBsPxrmL0uMzL0U9BEvQbYJ1DnK87nMQxpwn3GaQ6CujMkawlf2XTtT
YbZo268hu3hHvSCJZhUalFwdrrjQjvTiWE1mgMa0jU9UTzMsKShQPushv8xmGAxeBeNrSWrcU6/e
IjvasgbQoFmCLBsAZQaupJjqUzb14OgjQwe2Px3w7NoYIANi6GwRDYrIlF1a+yyX9pveylCEuwEn
SswdN/gCW+SOWvOcr+xVukHK7QYGAKQhkDJjRT0jT0oPr6U4QUpNSgUb+OlodE49PIOz1nTxupAu
hAwYj1B9R8Y/wA2fBz67JoZHoaiiYEflTOO5+vuAjRXicDF0y947Gb8KPQxnF4azhhINRD13Fj0B
64E27UmyIJ8X736AZ68aJS/C6p5pJH6gGqWhe9eR9Hfn/MFK+JVwVhJQxbiWkilqEdUN6oWiD6kR
LKxOaUREzDEhEG1y0+ZR+3lgEmxh5xR4XxCgbWxvxhO7NBV6jd/y3Zg447ShTjOq2bnf+lwfebbD
pdTbuJy61BDIXA3MkI6gM+f2GOwBSaCImJNaaGoQPEhRTdJqecdADGLKtyivlhoFqd+arilpSK6l
h44GTdmGHqPG/IAsYrE4RPERBW2e1b49pxxMjx+GA1kNskVz5udLEHUncVaqFhziCTkro814Hbnx
d5OxQddD6NCEvMcLffo/bxVavOWe0OLhebQPqSCFbqR9kBQw/0hcX/cctKmsHGEFz93k7CKWmcg4
2jinEjNu3+c2Jgytc3gpuIGo3HTZ14Mufgu8x01rEfcbmSq68nbc1fHJT+Jcm/jsr+nqpnzWb177
iqItzth7RSoYmWfYwpKw+ZCGGW1C+U7LWYX+Iia24ugyTGRrlojOI77cmtdJ36YVSO+RC2DykumD
dQFx/apFS/HMCD3g5N3zbn+p5FEXm5ImW7KssOW5ih/0GW7zNtKq9Y/65ExrOZMVjBE5p4P2vHuY
hzeQMww6BMWSAbiI7/ejz3L86noc5M8w8D4zAAaMDo4/rYvigW3lI3eVkOf4Y1RilebNjRO/I8vN
icJUyN5QGJSBoeSIJUYd/IxuRblKAJAP7KYuy+0JHtyaGZqu6EqMI9LHUgtBIO/6BAwq81HeAHyg
TGVB1FJ7obeSZj5VzhRdrUs+sIulHnmHgm2H2rN4JO4iqrzENFPV3gVxWA81+dEwCSIrpHRwSAki
KPFiaj0HTgNupSijB0bEJwxJh9r4yhlctZs6gdlIyPCt593XdiJcdkmCNXFeoJylT33w287XWaCh
5H5fpiM5rAYOfBXd7UbvnX/lkOkwks1o3MjJD/45cztPwRUcYKB/QpNO4MajkWniO1ig8jwRWIUc
gSD46RYKPIQoMZ7r3JyeYCic8WDOQurY4/wUMUfMTlyZRi2gPPqrJb0qZKGJ+XUL621Gg4RssdvD
3aJ+7NHu3KWaShiiAm+lPq1L65QYcOzAStMmNtGEClVgkvPDX3LCXjiZhecjP+l0MyMRqDQpjSL0
SYMQ89H8i1ewA4rjmyW6ARPpBcfH0ztm66HmPCaDDf6+bfwyFRnlHZeoFVax5DSs+EtfGBDWcfNm
WWDd9aRSqDW8IZrtKidwQMFqT2qqFBumzlzRYkAf0JmYItOh3IxaQ0WsR8tA+eUd2qHYX+xN0rIf
2aBwkPJ8HAA1Bw+YX4BCZ+ZfppCpB5lU6WJ1CT+zIyi3JqAeKRdNLb/wkb0nOvhFFYmHdYfdbsgi
2uzdvdtJunUr5/RfWaYgAXnKikMhk7zQWd6kJwtJ6pVuB83rxq7LBSzAjtKpeX7K5wLA2eaerkLI
plx0xnBaSS/N1LE0oolnSTbh2iTrfC+SkeEAUO8CYcSobwRd7d7HvMkhljA/OxzLriq3asxeRy53
HDY6buRa3cMCysyllBi3OtE8Eq0lgb2Ll47hzMG5Hr+hloP2QkAj44TGkQD0OnDya4LU1wJFgw4W
QM2ms9zPZXjg93fr+XUebi1fUeMa7kjlSH8zlEqZV7rU4Z1pmiwiDFeQ2HXRH0hf4d4FQqeQshtr
pY62g4w8UZlAyUtv3woEsF2kmQFfxfp+A9cISCKfrdIXnXvGantmFGPYB4txrDPPvwceQAoartqV
/udULCzOrIe9vQt5SZ6uwNLVo4/pApXo8PIX58Kxn48fhVX38JSCQqsuakFfTt2ENh1mLRGKVP9w
eqxM4InqOrvnQnTPktDYLf4xdqtzqzxtIIEbBxl3cx3lOQgbkSm1bcaSY0xg+7ioTuezJAS/F+w1
VcrL36KhLPISz1QhQHkthslgnBuWSPpPdU0sZPcZvYWPsnKcJzFJs0DHlKApaBw39Z/qHkz5Ml3G
9m3ZhajpWAcdfgfvttdBNk5B8TnWM+RmvKU6F1xHOaNR4Ia+EmxqKchT2YSIIhBPyqlZztaXLfS9
2SWnbliiuAqaVcWaSPmje1U2KiVXWZShgEvR1qp6Nx+H14OIi1wVQznU/HpgcD6aLVBin8wdohMf
e/jLaz2lVL8Kk2wFW2GRbTNVuX3CJbcChcDGIgqKKg6QLBvB4ZuF6znfkBQCFkmPt9D30cbgazbg
h9TYoh7wk7Z2uplDkMpibFIcLU9Ob7frdRud51VOF+pQ291gU34HOCuNp+0u5rPUSWXFFckR3YAD
2bLXOPdv23AuTANMdITo+Wi3dYGABZEz7F3OCkMMP8YcW/vXsPj8GQvKEca6YKru/WW/WxGcALWX
ebIAY5dg+q3ktpqD71lBI7V8KCUiRO0BsdMtkiGLk02VUMjdNqFbTyAzy7DV0KnTJqa17vvhffu2
K0k5TmYMo1ce4aUwyXBGi99x/NKaaHa2QYqe875SolVIos7AIP6nbxHbdXvUaKaU+V1YEGqCwRSn
if5XiAsWhTqqsHDpeYx+MaTVwfqD/IbfeEWljD5cGucpYJiHBQZt5NqPDb08qFKpdpG0m7+w+t/R
y+eOE0QL5pOnPyUeOATzrtwnYl1nRzWWjjs4rusHTzCmDL1qmP5pTePq5Kzci1BndmzzWNRsdtp9
uId4IyC5pvV70z0kpr5C2S2imeNHof0bH/vI36ez4lPmtMwI6rC4WxbvcKikrxBM0fSqHRl5kEV6
61MueD7p+NApvwVjXm+Kav4AW61mzmMK9P0JPCo0GIDfnwDN94AUbJfb5bxrLMXH7iWiv35iaYZn
VPwdQVNLXi5M9ZxVRFmBQfmW+RWCc7PkZXD8TNGcYYWnKthSrL+XMSQ2zTzSarMisNI3BrdMhVaG
Qq/IxoMcJdv/oe9H1GKd5pP5zxP9iOH49VtCD0ZPNhVov5r0jCTV2XQKDXbocaZA4+PJa5j0eHnY
6cLQcKf4r5N6U2h66wlSDpQKz9GzThiFdmpAi40Zt8n0xyYAOHiSR6b2nXu2wPte66bE52yZ+y7T
uA8nQ6wkkxtdYS3FTaZUu8ya3d7NLK2ykBzgK94O2OnACpIll1JJV/CFq5i0SmsDzZu0kEwxjEHU
Pm1A44n64tsfdym6hzd71Gtfr4xNiP7o/qRH/6VZD8IT7lcfPaaUbh/VKpoeCarRpHt9i+zMshca
2t1q0TdP1S5jZkVr2/y+KPeXtk0ouw8XlpIHVtCZSwLkpW2+qZik3KI+0+jzY0yksAlCi+gdwx3H
fUPMf3m7xmSO5uE4RVt4MgdNxP9pwAn3Qq9PlKLmncp+hVCst14m0ddBjJuCgPOdDyawtZeufYOA
Cno8tiEzIy1cUpegZSUkXrEcsg1N6TUGKrZq+/dq89qsqHWg8qqlTyYRtGCXbmCJeGgbAvHycimA
NRXTGaJu4/ZxSplPq5FIt18zOtx7K1+I52LnF4JauXMwHSo2qYJJZlItMcySPPPPYtkfgv5Ojq0G
Ru0iMt0Io+1kvozVayMx5EEi1aceonDjG2OAGfZa3ts+euqGGCq2HMgMbBE62s0UkMw1En7GrqAY
33R035+XzJ+M9Kib1XZWoTnQxd8jf+AE0tqck3KiHzLL03oCvvnoih73UQ28KMq8TeZO6JA61eXW
K3HQszGEH35i4TOBavIW/jmIXz2/Ff0GOw8ljlAk3EZLNk7XD2b5hmiI5ktZMwv/jFceEGsj7F9d
kmcZ9WySfkK/HtvVqyFFSOr43vhIDxXTsrokw5uoRS4hFDswPOdkPBVR59XOeXrSqaVAP80sOwmG
k7wkEE2i3vNILtjHzYK0Lf9CGcj2OFYGywh/b2CQ56cnDE0qLH9PAwQmxT6fswqWtZBxxuxYThKi
vD0UKeqffeo72rnfha7LXJCAKkNGCJjTwwfilJGr8wzXLPNC0n+p+tbp97nulXTFGY0dqga41QnF
ujCzdEEVT+aBQ3mSE8E/qEy/ZlNSfwfIaGpJDWX30DTUumX1iiCJ4rCzDZhYf3aeMlOxpd8/ifGT
aqaTpsFVxNwQ+jt5kj3I0NKki7SoSjC23HhSaHBpXMS39f9nANW28BRIw4Eykl5JhBwkb3mv8oEO
iY8jMAnsUdT5HoC4g/mbRkqNGMemb506GxUJQDQFHt2yW37875gqMPi3t2ebCm0rYsBVy+q1S4Bo
9HQ9sW937cXUOCHRObccz9Uk4w7fM3fgntVzTgkS/TlzepXKnTlCP4wO7N+eBKb+igtgItuhCWQG
LObfDV+5FspmVuTsQEblau/EURGJ9DOeBqlVWJoQeaqPs0icftBauWAmiNShvJ5l1xSKhdMSMhr7
HS+MBRjMuc9LGWX21tixtJcfVqPLEv/BJl3OeTcZreYahx8lBU3jgRBGP1dIsUk2C29PrYfHHGqM
lyKYmHeUo1gPcWA5aM4b8JYNxpaHbGoIo9Vma4JRB+Y5PNk6rl3tpIIQyS3sNY4k93qaRVgfHUPV
0xzYZKqMDLO2vhKWtrMvC9TN5q/2pehfDaCmRlqYrdqK0umtVZcFsndqJXYbh0ymzcPabmHZt2YF
S50n48lRYX72qGNUvdtxD6ZYVvPkbdEjtMnBCQ0pEZ/j/bgO4UW3laNeeFKIw2BNEpjNnvqmBPZu
+H9KoyXjBtQ/xrq3jm6G/F7Q0Tmhur1DqYtOOpbpwnVl/IpDrl47Y921btj5VEfMYx8eKhT/rszf
jtcdN+G1o+ooDDVBnVw/V9+3EierJlq4QnZ6ctrOVg8hCo5pxoBApnnTIxt5EmvmkNpF765ROSeC
GnhAB9XaXbhRTWICd3M7cAXFSCHaIGODyW3b4yno+eH/osNtwk+jSOCzgAkHa8lUwKCNJF+h1zCo
/r0spOd3mOW5ejxRKNURPLkayTocG3N3tQZaOzaMP7t6qL+2V7zgVJjydUgPLIhGjF+HJw9obYSx
miPsVSLAfnQjEqkqfplwMzFYXO07cvO/sk3P0eyxlsdhU9SOiNp8Oxm/yuECg/fZxrqUth1Gb2/q
2nuypmqzgCdjlgrSAjd3zSWfnkFhCtXun0pF1oQps+BXuxhwniQqppCTXcTQZw6I8HSMRzGMajIk
SuOcOLSwhqceCTzgdJ0roVFoRUyWQnyfISjkG38tx8e4NWX8aUXYIrkPnMnbz8H2TMIN7M+hINaA
LSB4aH3qHJSLf3bcoyIF8IZ+BTfxlx5QzSGOdrnEZkOkQhkD72KOCvOel7qU35NAKB85yGzypDMR
zpMd1jQqrQ3QSK4d9g7i1oXgyQ2zVZ3FYXe0DmsivsoQ/CVbeNmOjVFxeD7nOBLH8TtXv9FVdBnb
6L4s+lXQDc/l0mQ6ff+ntmTPnXQYNtYoW3B/0KoMhOd85CXLab0fkL/mdP1d0kjQIM4X7b6Bn0n8
GEb+rIm+sBewqLunMcvGmjL8wYj+VBLngw0k+YblMGUqGeszoQ3/7JM1eOkpqe3/RIvbeus3dUGh
Jef581ctpBESyGEd0X/3EAO6FABmwg6cdANIM85Sj+Min+TfxJhlnMGsPb55Z7ImTLmnuaX+RA11
KqkHzRuWChJqhCGkbwYIY867E9HO0utIXuKNblgaIPtnf7Qr4whbipsO2G/ocCmbj6GAhirLn6EF
U0xrFHFS7gXA/bjP77omAO40/gbY53nElwn+Qho6bXxoGZ89t//cfz1RnUNgKZdtTqvZxm92twCC
7MP7bz7RF3ij0Mfxsd83jJ1VNYRTXh/Y/vqRiFIt2EtHN9PtZJYHTDnb0q4accvcFSJFGJHc3gql
SDZCDokDNRrpweOyc/FS/xB1mS6g/xwxACevAUJ/MrjawLCf4Ii5lvvINvdnIeL/pD2bptuugHOD
+GQOUNJZvqvOD3eHi43gxlfPt92aHgtWHKsYxdV091zndQy3O8cDG6TuxVVHUbakbg8aY4BdP8A8
g9sTg20B53oNbs9Q3C/g/fnE9Yv0Ap1USy0itLtKRLU2uyipb4fioTnbyjLgEejR0tXpgcXXuXrx
D+72KXKat4CJEXtD+d3x2aQT5VVcQFZhn9ZxBp1ThEbHjfLBQxNfZ6wHoJ7pJ1dVV3q8wptXlufk
ynXeQCMtqDeq9cNIKjaVFWg95smCavia8d/16dMZ991hfNHHae0DtDCB2fQoc6v31ZSCmH1jaFx6
nG7fjvb8JkmR8v/COzyTBmwGDAIijD6bVvT8LHhpBYr6+hPy/A8JkAE3mmuDeK/TNwg7EgNOao+g
IO9y8Elll3uklmlyeWASglDKh4kdll4iY1EoP8POzEYvmG1VtHS//fEftGFO1YB9SzryMA9aeMXT
KrYg5MxY2cBGoHupvK9zUxGgxLgpVO12IYDGsfuzZJLd3ppPxrt7FpgBpQA28/SclwNfbCBN44mI
M1q43Y/Pco63awbROXThEFa2s6E6hLhDA6eNMjqP0dWlkWu+dYWbuy+ApKpkBe/NhZ+lAtSnr3hV
p82MjZpye1M9bgSjLHu4ZzRLGtiVdH0hp0GJM5/VvQA+jA5gYsvoUTrUv3HHOAs0MphzsBBH2xjm
pku2BsACyGpLLMDMrsyjXX2qy++4BqClk2M1NyxA8UV2xhdjkUKFtY2IrCWgBKdG5uzdFkDpmeVk
9tvnxAxp86U47GXrWVvKxpwAJhPB1M/2M5t9O68k1XVE8oh0/KQfmN4DaI7aeDaoyvlRWVoklNma
Nn+PWKsYgcU6YbZFMj34stjZ2xhHH6ilm+dOF6xNlVweaT4NfctjeRyxKdJ2tAkYoG0jsB3Sdx7r
Lb11HePh/PM2i/HVN9tfP6v5eJNpy0ZURCLwwsQ9o7Zt6ieiTq+MGjRXGuyJqaX1cPa10EvIGUnF
uB6e4ktOJKm1n7gBpMF7qEF6iCvlmDTtyUp94EyaGfVMW+CIiqDSeErnImc2rPk/DZmgJuuJ1HRQ
Z+nMBUJ0JS32YpJZNASZpL4KAsn3BzRVFLYQFs5hSJWx1h9flxVwExI3XuC4oA5O+gQ4zLs4qfRB
D1PAp6ZaN9WkeKDZebWk5Gzq/4AkrM0f7vHZ53cazXz38KTtBVbbs714QHZl45yrQjrhbiIabZ0B
094/gOlsRXt2FHhPvZjPzFgNseFApHnfqZOhGQ/iT84/X42RV1TflaIjOzt9/PSVB58eFRE3N60F
jRiFKBJUUm01Oc/q0lR6aDAubbuf6YQbltykVbVlU3GIw226t5TrnpRnKh0KZGCDiD/cOxpI1Lc8
dgln57C9l48RvUkKmweExbk1L+0l+t/kjN2sjiRD/aqMA8rBrRuc0ltR0zG9IWmm0vNzkPus7VlR
qG0qpYpEpNOLcX5dNRNbK6OxFgk5OOVUFyABeU4QUMiB+9ln+2cDYtpyiPLcJdsNfDBwKTi4Lybo
pdvR3fM6BTGbWJwqm3IfAf/m9HYyJZBYVTsGQJM/vHWs8/KpforT2m8iSB1fkQlJP8IXmWCOfjrT
qx0S+PSXVIqArEZIRDMAtH/+LXqli2tiYZ2eYYJDwjtn/3BI7K/rQbd5hu6PqxAhT9pOqnDoCVeV
gfIu5zp3DescBe4CG0HWjH6kW+sZxvMbYQbVfvezrp46rwcYusIDmvVZ6NO9cMBsy+IUitUTPifo
vDuwEoZj9VMwLdy5gmxUilY7Fr4ViiWwf1vuWR8WroUa5R3EnVKrP/HYtzWk3M7DhurTwKp92/fZ
ThXR+0+w/cc+Ma2/MYFbEpxXaNAyMcjRAQVSQU32ucqlNYT/6ykui3GC2IG7OmYxG1+ZTNWIyNNB
KKEQIB6pIDpyXRWe3ZJyqhmhKzyHlyqm/+PePjOwuBETH533uvJ6PAyPU1aqSyUK2rLXZ53XkyjX
LRNDMExo3b702Zc57SErRIEegAFufUVH/fMGuiDoQ+se91uy9W6jX5XFo/MFbkiVB4T9xtTTNZig
Pk3+S0iUX/9o0RZ+ltxr52Q3wtA+oV9ugem10N9kunDPaxEYmIFscqkTI867KS4l02FVHulhr2G0
3U+8npCFSs0mmn6JPNKvYormUHKA8yOFrVZCJgOG2VZ3mQ59a1IHFZ95FiXTToW6R6XUJa3TVNh1
DUvzAz8QjYd4tL8O45TN6kJwCCgvVbKec4P2puIrjF4J8M5POYZkUYyKZkbk6m/86POoy4n+5fBD
Pgr+iKeAE9xU7+zVgAE1BFcSSL4pITtewbh2ta9i4Wp7Sgs5IIHn9VhxNLud4XvFu2ruKFt3mEkO
VpDF7NOUUDhp9x9x5glfk7iI60bRWxeuuPQoiqbY5z+U7jSR5Pw71qkRt5VM08c/FxMpWp+1JgHh
NkdJeOJVAthbHU8QsXNbz8gk1+dXKalBucQA+s//y7ql6v/8IgRMHJVeJpB8U8me+yOtWzC53wvY
TcvmQGi2JOmmZ2tBbFWlQ1c0WR1ouyU/J1+gsIiF8a+LxS+gMjvqzeJNbc+BzW340L1Gx55/aIMI
k31UjKfwG6EAbmDasP3Xw0gdFqcIsGomprVWcbUNJIEkCQi8cLsdvzsFwkJzQpPvVpF/Wpwo0NPg
ZUYcLbyT9cXojztH7/yprtoWNKu6Y4hMAf/d4ATh6LTWna5gAcWP7Qju9GGk+w6+/1/iTkwsuWk8
UAwyMk83Vjrw75xaSyO8ZTJzyV/+w7rd4ElXF4pMhss4C0bGzkl+QwyxyZ9bhkOBAqcR3FERVB+/
XG5fzUoAyH+Y48CxLozjYriZOTa6gC1usCYPbqZ8epepULs6HJF7hVzGFtVytLbznMtAG0QRf+4s
T3xwclYvrmwjNySQAzGKydVcMUO9f3fjq0Nfm+pRg1qWzp3uhaY52YFPFYNhbvE82xh0FbDWFCQk
hyHletXmmv6Lu0fpH8iNfspzeo/rSmSe0Fer6qnO5YesW0ryESQ/mTDg4oQMq9H8r/7fwWt1D/qE
P6hIFYG578UlrKbukNwWcGRSOp8Jo5cJUlySeSRoSMRnYMYyVsySpfaOPD7a6ZFsxho5u9oIYFjt
b6oFpYKGL7+q0EwolzIs6qeu5KeZsdoBiMrdcKfUltTgWTAvhx22fJFe3JEjdAxJCluX/gujzF0L
uPYp0RrvTDpPpCYwuxAQYqYA55y7yI76Fgab55dEcP2s3hTfNeBIupRW1tJarTCa5qgR+BEXWtdX
BsTDI/6XdipkNQQ4U4r+LEBUFiJLVhSexVGTZY7L8dW9PxKpN/GPLugn8TCvK7P/jDFH9fGUXwYx
bTKpLnkFlTddy6ueLCDvt+FWXJIVsiSUgPp3WA8CHuGMxkxjP9IbYJSx3hs4LQiUzgeZtIBe/5yC
saDwnoAaVmJMSqbYs/4r4N1NE2QeUqI3U9xB3uBfnsg1Ew3XTBCSPWFj1X2j4jbiOng8eAVDnl6q
vKBJdRScs+MoZoTNSWGNpiafEkx89NyFHtuCTq/nNu8oexaOuW0CQOmQw6QnDf4fWc/XOzV51J0O
NsXkx0eI7HN4QpaW2cGYMwybaIvv4jxAJ+7oWmPHgkg2z7QnxbFWd25Ggo1oeLdkEGI/n18BsD1n
664kbHjBUcnwG8ukYemTYUYSHNUW4FJ1hIjAwZj4kUvQgMMlLr0BwtH5I1pdlUndNMyA/2rHs7lD
AxwpjvqFTrtd+zvSoRmn2gYMXerJjA5rJKYbS5Jqps/P4bE7g9pkGYbbFDbjZsYvo1cwepIfYLK+
ijttrc5NKTqUmtP4DYVxDpEYkX4zxQ70NpF5PQsIQLsUBbuiN7OF81UVM33jzFraVXGjiOiOxFXq
7p0cv+L/9DauvPQ/sex9u3ae7yooJQXUguGfabgCWOoqWvwWNDD2sE5KxV19bCtDEyAJSoJTRNwW
yOwFVej99BzUeQDzI5lE1SXGiFBmsZrATS6XSBadTZ70ahYgVmEqKDJrACljAyYg6CtibgY7xUkd
NzMZ9Jz0Z3DRWFZ6zRmnjCZa40cPCmx8XeiQzO2T5X/SF99jTNKYFs1Q7L1OeoEm4KCgKJIp+pc6
MIMgs11AF60xk9Ol02r7bvtP6TK2CvhXqNWL4oA+/0Gt7zOHej/fv5vjYlI9DXLk6Y2R1LEfUigf
tpqBhPn6YNdg3L5J0fd4Q+oUui6VGR5SZJTcMKfopR37SgCjKqUi9vBu3Cs11HQK3scC+hscqkXy
GSpQbQtA0/GFWh5HOZ3YyE7V1UhlD6fVapjt03uThsRyY7u1gxa0UUuQPZ+qv5QEYmzS+edH/bDH
O/y0N+hbcN4M2wjKl+TAhX8hz3NGCp63VT9MxH/DVN+PKKiEBlm/a0ryy3hXyMt3BOKH7r26yO18
vHkMTn+uAbqsgnhoLu3iH1n4NAr0/gFjX2c+NRDqrAlrfmk0u2NU3XXYqFJLIbTmnMRUytnIbZkV
4ln9/Zsty5ngSP2BJ2dOmUDMXSnc726owTltcHoKAvNfNRWc+p3bgfFvwTcs8W+G15jqum/nsCtA
RhvCaxTIGVFGECe2u5oqjyMrU3x9lotWeM7QNv4tSq6TJohxuPjr3PbxHx+6oWl7e6d3UQf9eOHZ
9tRkRFjW9SgknfZ/rHZOjTZBSw8DK/4cgbaMLYHXPOkvfgZfWaHuFr99K2ZdO7cNkBK+j8UDaKB6
ZIRhzwkUW8L4M3tpHvCeMUUortI4bGhq3Zf7a9//wwcSurPeE9qx/nMHPaWJ7n+cxFBcCDboansa
ESwt7JrXpPeervWq/cQ7NMIr2wSXumGz9oH9EHYkGnMmIx7J84ZZNnEeL9gV/WIH+IrVIx2oZXxc
/XON/hdnsPYieYzcD2W/sVDhdA66E90WqNf7R2EW2MlW2Vv7TA2AY+TTtOc1uyHLHbZCCok1/7GN
kHzH0gBHQ90tUjbKYAXj0X9Eirokn6g+F/SNmpfVlFbdVprItFKWSF9d3n7wvjC5SWmq807C1PaU
ITLp5AV0LUbcCKZZe8m/nC7Yd97dUOOpPgK/Plrb+5emewDVyFTwWJDIzJKtd5QNoWBWnxhUf6MQ
kKMXzAsSgV8+rRqEXytRBZ2Kg3extcfj0uUrlXkH57Q4ZiKeQic0MVkD7c1nY1U+sKfDkMK4Osip
X0mbpYbWT/lsKksI0wJ9TJ0pHdsN+CObAimVPBUtWBZZ7Y+fivPG+FkiBSmXSL6zaIEe18scfnIg
NNqf28h5hWq2G7/lZ+Uxcx1fjLi0ifvr+ASJamlakTFTcvofSFANPjQsmhkLghZOv74QfrWTmalE
xqm8X2FD1U08fF0P52dqxvnbzUUN70u+cW3VTSRsuRYh/Su/JwbR/t3/d29+bmU9z5cUSKHw5AHp
iV/E9HDUeuKLB94kK4c1cS2bavNMIsDUTHOjpNsGMTT0MPuzSmWEv6ZcAMfAc+Y15dmGayLMiZi1
SFvpbhky1+E+WBhFzG/Z/bRU/fPF3autdBrM9cHY4UpQ+4ljiFCD8lTbztXU7IUILRfdM3md2HrY
UDceL+wTjJD9bcqDQKN0Ukwapm7SM2DLpZw+1ZxIREbfl8MZGppsvVG++1gDQPea21FfZrV8JktH
CaSROwfVkwfn1pWBuYD6sXsoqBKapJZcTdjUvhZl2BEG6MXhN59iiDy4WLnveB+oOgpoWgFY2PQt
DON47diN8FlevcOHQByQwPFbnsqjY51Cr0rhrAvv8a1ytll9RRE6x9xu5pmOTZF4CSe9xi4ljY78
yPf9FpYJLcIBBamU8DFJrn5X+x99+ODxT1FARFkK9to3R89QSqt40horCSQRPF/15mCiYB5Ejcvj
Lkv3ddBFph8LARDglClGiMyqT0QRmVe1TAYHnkJMdpLjw2Ui+/GEwTH9BNtW7WlEgPtLR5SDcmRp
0tccFAd4DOgEpXiQjFUg8qugqhLW2aTd8o6Xe7PqSxUjwUOH4MiVO/XhZnRqugWd8SZiOQAdN0D2
576B8M4r3WJbIITj3GZVW/bSAwu7CehhryfchIpMR1vs+8Z5qOAJsly/pj3GfcBXNSjp003+/BT7
iLT7MdLGJptm9SOkCrTAZqrURQ3+F5TSnB2da3g1CWQgJyNsAMI1o651q8SZ3abk2zRmAyUtL3en
V/laxO6ZtM6aoWH/NhO9zYtxEzOAws6dmilcA2Be5z3bemQzm/DROeTIy3b9lsu+06E+wP+euohR
ZSAjpNG8d85y02PST6bBmou39WWw9G1Ab7nqPXCK1Beq7zIYz0Bv3ip4z8B5skcTMCJZP7ttToTk
RJ9i7/0zG4IJ2AIXhR9ruvVZOK0gPOJ+T0fCmNKipNWn5B9RvEjMNLBKRCWHkT9gb0G8Q6vU0hK3
Vpwqqbb3PWwEv9FIgmFgwmrtXrajxmm3wt/1tUHpu0ZM2AMqR4rpDgHh+NCQYGveAVRMmZRELYOO
FLXBkyIJtw+VRK2gMHuU2t9WhCNqpdRnx5NrTinby6K3K0hUp7gaBB1WFXBJHSRLNVnrnFwWjKxe
gf6DrKiNt363NqzOFOz3grY9qa8kQbnShvk0bnYqxfjlyNpvtZkD2bnpIDjNDM7wXG1pgO8jDbUF
DP9umG2y+qN5ZvNZDSCMqntg0WTkhSKcYkB8VeiZTvmixaiNpY1FABl+Tf/8yomf4OPJ96SMVa9v
xaTon+i+D24txdVGIAC7rgVkCpikVbyP2sU0oLFHFobmrYCrhQgZUTiwKZBJ9vAHNMyqbdxM9Pby
apBwqMg2yIT0huEpkMXfCyP/0xDgxNrk2zUmIjNNXtJBI3QddoMnZ7utX0UyvTY7xTiT1bNgbloc
JwqP7Mipx9J+5YXtrwNQtvvj5XKZCYAewqJG5XrXQZwgAdKdWqSKfH6nn1azUEpMoZuZ1HVs9KIc
ufWfuQOyXqCVK5R8IC9kNSlaI9tbGsbDnW+GBXg37GstSh/qyuRMy+lmjYPLHi+3rcj1/QGFLSk1
llSH8KBLjm5uRDKuZ9d2TVL9SvewpKTPz57nUu6lATkVTyh5KkN7IPN/dUb3IArQC1S76Yv0UdJ1
mE5btqO8CTNqjfgTAo7utDQsF2W19R5MDAPYCYYO35V+j+u8q6jA4CyWkFfBCOgc/Rrt3jhxBqaM
73Rv0C3TpyM/+sWlndhoOonS9M+f4Akm1gBKXeWXMBdYRfduxqOmTMnfUBH+39QXCNw33/FoEp6D
RBURQ/U8CHmDFSvBxene9SgYT2ZwJ8bQtHr9W1QcWcdFy3oQOQZ2ZJCFNvl1EJHcyjZVisflkGzR
kK+UP4O5zfgBWOOzIJ09ZmXQVBxubsAhmDZVX75V2d2te4T3vSkjyV7Tx01DMVXiY2j0iRR8MoAE
lgnJ4IkvDnvE2+zQ01D3jhgcmHjtCVI+p9mBhc3wDW64WEoaHQW/JZ/idJ70nYDqPdMk4+RZiK1d
qko+Wa9LeMx2HsaAFJ/KImXN6A2uIr80v05gLFTgfLRFodyNk0FGhzwvdhfHWOc0ox+WMY3y9AoY
bCxDS8YlcciwmssHqCoGg96fSAhObPl7WUHq98Mxw/irAl8VIx6aqrYIBA7z2Hf7g9rAayglJVB9
v3e7G5fFLtGKNbOpH+3OIY3D2U00Rjs0AIBn48dsSQbzi+AS8Pa6wYmexS8Qr5XKBqAu5jOCPEi7
T1/cD4zTzqZ+8lFtCYYPVaUE5WLlKJRvBukPK/6+6sF03hHiY84fbLW1uvPkd8RpUaicCG8WKzyK
tDhoI+SOa4Z1m6HPHNsmqo9iUTjnqqpLBpFdtilkE5rORgGOoC0m0MabjyTAuu/VOHjehv3pFbpq
mh1jJW8T9VeXifSomw4+kLVYUbeajm30vPS3zi4rqLymfwOcEpXOv8fjMCOgwq4iMYLHp2JQUf7a
24njOodSo39KGA8ZdCHr3sAivPN6oW05nDUPhp/FSpcAko3+h0qH6GneXn1sHhHYnSaz6DB1xaKU
UZ8Gg1GcnWQ/5uaOrcY6AVPu6y0YVeQpRDaNUdR5HPOZcIJhQNna4Ju9nu61goMDSxWBwBPRJg/2
n04tj3PLgyFd9mBWt0plw0QERZPSC5QkUcLzPNP60KMujJd20v5CwRWMazULUyczCisqOiJSHoHG
LCe1OtcTfkbszsZkUqhgqueNe4aWeNzZGxClwQEHoWmMUFV62gC6Zaea5QO6MuQx+4u45geUDFaU
TqWTksod8JpCJM9VhtWGU9OM36JIiJc9Mv78WpUqx05NPECtZhFExdwrhr+rK0z/BgW89rDvi3C5
tcQQlFHKs49vJyvg4krnUHhll57A2dFrUSv4TXtX0GDN4oIjG21QzobHF+EObxqrlvaJrtbHdheO
ybpH5jGw75gxJIEjC0cemU1B8Sgk5AtVBIWCVCnJWF2gNloWYkHV/1lmgrzWfDK0FMa9tVmmsdZK
T4OiQQDEEuhqgSZI76+MTtcaSbKVOtj6DkfDk1Tyz9LdaQAVKsjgg0krXXisdqchIWiIxyi7SpWs
SSSufgDItGMJ5EcGWwPlup0Hope6GI8gyWwxr2MzR9I+whXuCCe6Nzd4wjfQ9LgSFgj2y9kMfH5T
+IksqPlWogEbfA11nzI2VW9SS1VA40hJTVFl0L1KoTH1oSMgIBvFQcqHDdSj4JHkPyW1CRoqlRmh
T6FXKHcRU/f7bbXu2DV7dUHdhA0LKe1WWMWSGjOwuAyfTTt/D+yOS9Ud3NPG5jbrRgdYvSRjA/N3
2BcqYkede4gIK5ZXzA3zV7ngJMs5jbkh6kkcGGLgwINr2TPuvyJlGymRS1DPuwITc11BHyOHgNaV
WsN7RoifCROIADvH7vNjCM5jpvwA2IjtHLAfToT+F6cMhVf49EXI3TowG3PTvPucOZrg3sfhkMu8
TzbyLsvVtmt2kKi1Er0bAdWgoJK3OW5/6GR4Nys9sv9nKLvClNWMdhy4uNIrq40JPpz7pPB59IdA
SGVzmlFb/Rpmj1dXiaVcn+cLl3cCpNMpFKfai6G/DrR5v/aBUtTy5RldWgyjVqWhzfrdDe1ve54n
xo2MyrSdLXi+YNmccb/foSW8W9Wn/Y/6iyMC2LVEFT5CzqXeOqDZbtSVe1x1IhTzaO9y0nz0ouRY
bZqyciBBds4DqCBcPW3jWZK3ZP7uVzxNlBnvn0snod9fwcMNoRrCz7CsfZpmsTUy0Loux4h7uFKL
VtUK1zw64xAk6kUoVOaYnbNuzMnRK7AV0QLn7A17t7sSQUbxD8zIvRvnQXySTXQ+yxsnLSe0SP2D
rDFInxwv70sJs41lcZjlIkfELaFNXqWcGo/s/MmbK6MrORet3IcsqZiAhRj2M5lXWOpyoYCMkmua
a4LSNM2+dTlJ++lDXZr/bfMSeGxyyv95HBB2YeNVxHbxRYOECszuLrldU0tZ1sKuuX6RkDMWbWZa
6S7qCH3HfsiSQBZDrwRtHjnd3puQYgsDLUFwqkj4BFHUexVqLFa3wl7l25ZUKs/CGA/hpSOujQc1
Oh0/oLwZnn/HXMEu1cqaj3UnZLgszpoKektaYJV88TrUKMVVkZfyJwZx+OFWbxGPM2ZjxTfGSwzh
aEXZluU3rAkop9frJ87vypDpWVxn3A6qtQLQl7nKJ841sku1kf6cwzYnLjpUBMhO3+IdUa0YX0+H
Si5FkGbwJenl7WqEJD64BBBSdSr0r+sRHZW3ZiVbPO60JInBaLvYB2qsa4ur7fF/x5ulYHQlOF5v
ctK96QbQkmMrvmlkpitCoVFHcIzRhMWZVrQD/LyzeCnWFN3Ocxr64S/Tnb7EGsN2NcZId3YsyEBJ
uXjKg7vRdN2KLOqzZ9uSNTIa+h6+fnJ3rSw+S8z1CIzgICoAVeT/vX0fAxQ5SC/MPIrdTDz/UkjY
wIewo3fs8zkaPRtIuEBhSF9zGwBtWSr4vtVmjUAm97v+7IrOa2Ejy1jzjDqvotUVSQb0DUfVQTFw
HCUAZK+znv+CzJ3ppptBS1XRHxK477MkN/rF6+YSErzrf4yBxkX7o6rwxFINUzpQeLL1/fHj3oSP
JVfF817yCHIRtfre/UJXRk3s+7V4tR92bN/nTz6Ax8Oo6ZKHoXAbTn4FssPvoTHDl8xJxlWygKUp
m/0+f11Oh5Z/4q+u7QPNvK6GvdaYdZ9M+VWRivoOFuWy1q/YjgsnFMAT0smC3CA+8hiNvvn87S7Y
fX8tiCetnXi5ODI+p0UVoKrp+uLLJObZF9bV85UDib+F7drpkl9MlhISrvf7cZrldN9R5S3QPlsm
ecWYwDSt2aYdK72DI7TpNd7Af3wHcaa98xv3tSZArNipEabCB+Q+UAroVRfHqsx5FkS7mmRgtK17
YBbON//8vQOuRDNKXWa1wA0EXEYzhyBwfRP2KDAvTuQf2vZEb0jAixyaXlDfDiZQDmg/Eri7S4F4
B5yeComdhZRH9myyB+foIC+vipoCqZMvaSfsui5EryNPY8QOni9qnjfx161RMNSb4LNjvAphq0VK
HksAnafXLz5GN+b17fNb60vboxbwf9m9XrN4mT9rzRycO3Xc9aZc6zqVxjGwx91OetHYbcv2nMxM
BQe/Ss87GAnNHMu0dYJ/FNyVK7Z8FNYX/BOULXcEZLHrWpO7DZ0rxBqfJYBzXn+/OVEIejY3h0vC
60rzShJEzN1jz8PvmvWuHQZF5LUbeLA+EyDvVrQq2kLTgkzYlNNtQShSy7jINHTuuiZKUhjftbdn
OEUKaP6mQuIJS8vVUASseSrX+SMxZOxWhnyrmcwyeSAVX8b50Wo5iu20DgVWvVQNe2QKcm6odwFm
VuTiHzLvvO1zL4jTguYR/dq9OMTwb3mma/+4Q8oBUjgPxfrHu2h6C7EURrKWkqARKZqfP0TIh8dF
ljaT6dXe1mJQw2+RRxYJd6JioobaQbIgU6bLNUKlUCOUT0W7InlPYwyHCjUz28rlaAgzyOi6/KRg
4mK3PsQhBtaiqG8yXzqjVNdN7e/UkalKDSt87UVlMZjhRwRzd8qukJyY+HYtmg6Pfff1h0nshD4Y
LFauTnMAoTSEW9Q2S6kzz2grTVUeOykGLdiLUyH9DuFxgBENOP2EJgaUfxoAv8qs7jeAyJCtgWL8
TpCUElC+CkS5CuLnlfIvaG3iufVWK3IClM8nQNx1Jfq/euohoMemVrjXAxOn7MIWIJIorTERP1rC
sQVg9IHJ8hwBx7oEhOcvxMgTP72ClNj881DoeS9sLdIsOaKf+9QbIGlSKIkOUDaUr8EqJN4tkJ/Z
1QgIM2XgyBivAeh7fnUc/qzHip2HrKor0KSQq4Io5BwqPhCHnrdHXqXyg55aD0jvgSC8vxz7tY1q
Xj8lQ0tuObn6qdKhWBXOCFqKOHPOz0BWBN8s1LulhEmMpDew4jsKnyyAfUAAL8aWMbouiJ4J/U0h
Ew+VBCzRJpNyzU1EHW5x6eF4o+oRx40g53uNAmSwFVXGkStBhBtPaKbDIZyyVjvf3pzq+Mnjm/Qn
2IW4OeRAh2dWWbl1vUxq2vzb4LKoz7cQF6YdXNydXJ1UYety+QFzX3OxWjc+9ZKzLWV/fsfqNjVi
hzDQRCRfMzs/nQk0a/I7nKg9cE2YO0bYvpZC4sdpQmwvT2xto17WbdleLUgC/uRPWlVACSvWJ6r1
T5oPmPfApSrMb1mvoBzmGkVGT6BqsPua3hF6ss9Lpo+wLaLwiPFBxkE6Gm28khulUzAlDXiXRO5n
hhn/CTCZFlkiSA/7a1+jAvWEHmAx2LsrwlK966OZgyQXQhcvlvNWyLX3+JsBXVGZ+t+Um2eQumIg
DdSxxFzNHhwpPfA1O042I2I9CFL0lZiy/rZMpatgLYpmukmqA5TujNu4Bj9YsABuZH/DAKqLVm3W
7V1cuLdXkZsTmQ/ItUcJ1UMVDRJCjPB864DJLNNeilNDbcxw2X0oTBUUrG+Y+TxuUzraWnIlxBN9
R7LApdjz+dhRaNftGeBTOgx1FzUnvZchcReKENIL2xQPJ4mRMTBSukkrRKldqSr9yH/fb3e4NLvY
tpoKiUS4x1ndeNAD7szkIvBgkwecu5q7AfJ0UXQT81eqAhC3/7dODUFTerGCYQ7GH/D7MCkBS2pY
pjRxi+D7PJSZwxGJ4rVMr3kMJGrKqwsWSgsaPMolrlbr0Mn3GhVdwzY3b0cgyztP2cVKjsOXJbEB
g8FlsYLddsaEfZ1iT7FRDwsM5ERkblA/mck6p2oG/zLeKJgDaFQZYMQwHrBLgrmayH5QW29ojGZf
F4X8Z0fZjxT1ABA5eCvL0ld7cwxQQRSR4ELe675h03Y3ST7+b7UAtTK3plXFg859ZALx6uv3plcU
UpI3U8NeUn/YkddlwUXtyjZtR9rq05eR3d+idBCutLjE2xYjAl/XfqxyCYnp9OyDmm7BINnZlGlR
oFp+7TDZ2FHilK3fJvM8zWj6ga3zVoKvwFDlI2Yaq2jHK7lmMh8lJFerKi/N/9Q/p2vp//KFID2N
Zhnr9rcgrPsuT6T748sS6ZeWIWqCuE5fhM5Sbnv4a52XbhPd01p7MHTiVS0NUr69ptvL1dmPwCCI
DdY0D6gEip0/NVC/NiKRgnat/vLKiXWWTWCRiO00EetQmTT2m2X4gkSAaLm5nR7N8d/ADn8x0EYC
f9BOcT1RmEGZ6PXe8hPM2WNLlDWhhlSTXWkqWXkVexeV0zdvwQKkXCQtV1iaRbWVNte41Zz4SE5c
RCBLQY8yFebf2mVbQzYklys9n0AxlfOnuLD0O7ihB1/YyXUgxtkVL4KTS9Bmg5sxiz5+Ital9tLd
i8r5ur3cJwt1ep1SE8Rwy8Dbr0jRTylM82rg/KbN/Mx3UMx9vimlBIVTNkLxETNj8zy53DydYzDJ
qsLkF2UGNg9vc5F48mzflIYbd2+SHcfvn90JQ7/1SwAUI2yqN6aYRxO/jZHJgMsOQlse5nfXoGFs
lB+CL7xvGtUYAV1Ct1Nn0xfR9T4THtZ6Nom4ABhLnNRY3I+9KinLm2m41AKtmpFMfgbVPvhLrNmK
GhCx9FrKHS81HWYnz1EzUc+J9eHnnDCSBa5rmRmJB5sFP2RXIXjEQ37WRdrAZhaNyC0ikEBNS+7d
pJ5C0mbYEq0v3jODckRcBv0PqNaixARUBvev0g4QOxP4J3eQ+8vlRJkee2W86RpVJa5J4R5r7ZoB
ol3koMyoApEjL9Gboz2HMYBZV9o2GZHSOfHRQxPsVyftyGiraw44wPBCP9K7JtezG0e6Z86Ufmtw
CvzIyJ0ByW2f6zK8aen8wnzgmM+wh0VEy/ZFXS/qppm5J6/J9xZgUznR/xCTnJvWtz+kpa5NSS4A
ApqXrUPxgd4G4AGVmq/VUDEVBTFFkObjhdQ+iwB475NK9Trojej6fAjwT1j6+YLXXTNCG3SI+Djl
MmA1sK54hxKJoSDTbnUhRgG+FkczujeuMD227+6poOyvCa0oPut8tYy9UsNqIMTdtFm48Gs44dFT
2xKudylSMNXSry1WTAx+0SgM7HKNG2JKvsptaqp4tINParO8e0h812weZDPvGZSPy2+qsU0ro7iK
dekoJCDiQTiu7Th0Nh4Lj9CpOmlISo5MSPobDHAPu4rVbSX0MjeuDGm2v/V7OafzGXNekSQvHy0U
n0YO0KxqMlyglaK4p31kM1MY6c4AgwWje9jls1FEEwEc9UxLf//g55TKiuVCYC7+MkVf0NF60EcQ
aTMCsoA2cAhCAt16+E92T1oRsbTzOtPpAb2sp35osKx3/1XnHn8LnOn5PL5/HfIsON0xr2PzfWXy
GNnI1eJK+N7QDS342Q0jAfRGyzT3ir+Pj4t/vPxxfxxM6a4FGZlOh81hYoilzoPfNDBNDzh3LF4E
KcNz5OdfxVdHJc8H1c4y7S62aNrRz6CvW9dxX3Z/yGcyiunA8rpbOVdutY7wSq6ikakUM/ycrYtV
lPZlNRTUmL3yIP/FvQgXqcg6vB9MUCHCpMqVBvxrF1EyC5AMhaHttam2+oKtltQv9OgdipwTdc4P
tZTReDX1XxWxug8Qlhri2SylZzK5Ili6fnDBBg+efIkSOCTF+WHQb19AFbTIgEI/t1QeGZBviedw
buptsu8hfBpmeinYzb61gDAXWz//JDeEnpaDCd+2FRT9Pl0c/oatUc6kj/xUW2My7Jfj4vaorvs5
2oOcC+ORdSnR1jN+uirASXJ5WwvigGYOkZbFeq+V4hNPD6spKNMHWyvg+1aUd538hcpbHHsSal2I
ekgm1WDgIj6eiudi0QnXkrhBQvqNxtV222d0gfrtJc13hvxpEjC4UcqcjPl5g1k8sP1DTZ6Vp6xz
MKcrHPqyAa+SiN0mUzaHF5KZAklEMo3vMXiV8tyFd+vEcxR+bf58rtLICYBzBDXZQvCUm+BsRyq8
v7zVmseWflUbOotgMAOcecWJebifbPf0sipQMEgtG0EzCguFrNnJEsaVLYYoTkWSCggT8eKvAkKE
rsbEYK9+AVhCyUWUlf2H/rmrOaWk7bMwL1//ZA6vQfuroSESIVBo1nGbiXNtNAlecbciPsiQaVjb
GoBaZqA4wt3UmeBAI6pWsbKFRs62b8WBwmHEC2Cd4SJDzqP194BGOsEghJg8HE9/O7vrv4AUOEJD
8++gZzuroYio5sgsrlPV5w/ZAMAqdDdOXUGPmscTiY6Xh4yRJNhiZia/WvUPNDADHkQJA4ZJZXk1
ryBlSYRpyM7/VDQIIMKoiUKckBf+zMkG7FqNidwo37wgFPnPatejrQmcIdrNmVPQg4YGNFPJ5yMG
Bd4O0haXu7vkltqSbSnLf1eRd8JLU4sFCbas/mbwvIKrJE4P+3Wp1t9ZiV2uWQYIGDpqnfp/2tcD
ZHZmykRyYlqHsiMZ5jYi0Qo86QczojEJBfsVi/ta1mZUNgdeKUF6H9kwdMCOd0zmidmN97NjA5pg
PouAfq77eg5W0J6pCs5xqeohopsqv92Cvy4+ReLW+5XNtoXCVYmvK62bMGeNLYLMG+q/MY8cAaXM
jkv8jZ7XI51IvMD8ixM9ymYARuiDsaFv2J186EF6TNUoGth793REUnoumSYwlXPjYEUmdZ8NdXFx
iUczQ0Wm1FwbJ/GrWZZY9pCoOj9oOM4BB0u8UEQrLONzfZEjuYKiNZ7PkoB0qaa3FkCg2q85/HHk
rP2EGQbo4EHP4DggG/9BajV7v5LXR5Dtal2ypSgqttDqWLG4mYMRAjKESscwsEKff5hAqwuQwu4W
9/Fis8W4ybF6pafBiOCOIunzrBoHHT4dc75cjIrIpMzzGDJFI1RkcrfAtJ+aaP/oL6iWxN2Lui9N
uZxS+S/U06iTlV/vLNhPdbMQTIJOyclEl6NPOBWNJCooOc0epUbpncK2VK43k/GJQGeH2O3zASJO
kymSxkeLLo922kd0R1FGAMMnUa+rWus4TqjTBLqNTyINBUdL7lgT4ijMp/FgHo8V089hnJ1EKfA5
1MjVjNrkO6tUPuX1DGFx3sJidrZdI2DWkJoHIc7k3Gu2rp8WvfJxiX28IEy8RkABfonlUqpn6fT6
7IG7fUeUe5aDnTgAvyXGprgSMxCxca1Jrhs1FnXL10LTNw9dD8J6dhg65oJboPISuwH3tw2Ec0+T
MECwzbJk8WGdDhX9h83rHeKdofIlC/yLr6uXwY9bEoF9+W83TiGSjNJQsJtQGKXExVoVONGcpqjp
ZfZk75QPH2SWxuR0rQeY3z/hpbq9XQnPYNNCXM5QPFbsVP+IHajrCwxPscuZfStzIuxQPbEs0ioC
2GOVxwAXugrYoJHpubqCrZygEQmrQ5mnnSjoFgoqhguFt5RBcKwZqWkj5pwvqpshpGlPnynViAL+
q9uRdaYoIgwXR/P8R1M1UO+zz56KVJASrIivutHyrN60TmUzqN0ALsroHhLPdIyEDExmnJCz1Q0D
vijbtaGhmOwbAaNiRDxT9tcQI7KMalFtirijvLqc91wFWDcRnbqQ/E94CiZ8C9g9moNXOeGWrfk4
X3gIcfrehUGyk7YxTjfZoS3kw097UcQ0OQ7MnPiiPQr0V01wkFA7rTSzJyCmka2vQh925fa7H8yf
ToM7pStiVDGx7iYM5Rax76YFQL4ICMejikU4yykbLxOWGc++PzjFUL2eRlP4wubZkFnfzOUAKcA2
vqrzjif7FfNhiNXehwq6OEfPZlhqjxNV6hGn7WkeH0c+bLVi3PZZcshrdSWhUhrhhnChyiO1TvmC
d7spph8O7Ep6oX9yCPvX4EgU54B6l7JI/ne6wlFSe70gdrckCSSyAUqE1OgkZhNt3UP6uRT6JXJt
W3veUYQtOcPqnUgyCFR5fcKqb+wjYa7I1TytWrhnfDo5JljTVCYOPFJds35dTNHPVxDlfmNv3viD
wMiP8j3G8uo3TFRsIquZ2cnvT6c1+WurIBF/LfKhioKG05uNLu547ThJJz++9BpKA6FeGe/eo6It
WHtjZgHj9f6UD1fKwwtt+bFd01/t97wNI4Zvci7w3Un2Qa8RvB77Ar9r0n45E9IfWZKiL4rOXkuA
GtUCTg4WW1eGasmndtGD1e2VX2uGTmVNkH3HALXpzIM4JMkg+xGVS7Zkiwn9c04SlLFf375O8cM3
BKrEm4Z+RJaZlp+zee1SePq6n2OIKvJYBiau7F4V1em+A/y4d/oeQ11ODBZEQTMMPDjVvbHyQbAW
dhEPiGUqONgRC75dNEN+G3m3rENqU58brvG/3K5L3f+tfU4rXN9HXPHTHIX/dFJH5RTrJxb3JTjx
WL4+f0ve6mH8eyK46sZRMJEt/ZSVSuzIh5vLKvif90DskeJC4zkblreG/9P7G2485WCYggeDTLYY
IAE7hBBtZ2Yy2kO1AYjsqDGMSQ+vtp+VPum9zi1/kBMuu1WF5k0hH3QNf+V5AjEwo1GJfEq+hYn8
vW4Zh8vzQaVpOEyMp8BElVH+V9HbOcM62bSeyM+L2CCul6/TT7CmBEtqYis9Nv+842TIcdQwjfxS
GR3vABihuBLgG8jWXdevz02ytng0Y5xK4hwfRLHVjVYj2WA6SW3nsBi+ee+oGpEeUabe54uHeHEs
2zpSCTLI1VE4UUmmZrxRIw6RT3YouuULGeyRelQu+tyGnxHgnjC/5WueLeXPJrzPf+pRSV1CZTjS
ZZAj++/TtYe1CZjWmqQ0XMoBFokdp3QRtP2hLy1XZuffMut1kw0dvD4gFT3YwZqR5kpGFADtRFwY
V1QyzdfTcgA101GkMjLKJqWDT+Nw5jI7Uf1+lzIlX67qg4foltGmhp1dU9mEmry7s2pI/npKR1ug
FQwmUEe25HQmi0gkCk8ytUEE2XS7SFGPO5pl40R2ARjHw8PUEVXgBKcaywjBhGseipY94mtInuKZ
6Fk/dVu8FvbofSJ1ERzvbSq8OO+d3OXvloWzNS3HxASgqc5UNt4kADwRLZFLVP/ouo8+SgCLml8J
PnoVGURkfo4WuVZfUWd/oaU73sNVaV/EA6+lj4JdCLjgF2pAER+GDT8ba/kdYYZ43lj0AbqjadeO
tVDnWcSyBOugwg2+xIUKozQZSgwtszsnjcwCDjTCTssXXYpl9V/P3MSVRLNPifppyH8VdD9n1YdL
1JfpDozMjKx0+66YrhcbNXmunOp2raXh8P3Q61fzOG6AliTuI2HcFQY3+5Z317tEWO8Q1tuB+XxY
o5NlsU8Jf+M7Uiih6ibAoHOQXUdcuRisz0cXCTR7+aifCingsvPe8gguZ+vW2Hdfa3HN5LF5ofoU
bfHxT+/kYjZC65hDMWx8Jiv54Wsp8EzPzbEAPNNmFZ+Qp+DTS2RF4AwKLeZjAQp4wFePfKgtjS2/
d76dBeY91o7eplZAoBI+lNHhOCMu+rrK3FPPaNe3jxs9rHyd7YlZIzhBIR6SFtVy1DvKKT56oQbF
VVl6UoOmSqpfTnt7rtskpKWbg56qvvgUBndAyBpRQM0FVGmKGM8ZrlYsw3Pw7iHtwKtN3kL5/65L
EXfTPOqPdfaiZKjO0Qe7n9mfBYr96I8HyZPhdyay65Eydgvq0f+Llc/TWUU1BotYdOC0ADNL905z
/6gWwJ//89gkFEICzsQwlGsFvOwQrha9DoFZXVQxM8s4B69ePppugKI5r9J6U6lcGeKghuc8xBoe
Prq2D27VluOYlia3Z3q6mtw2qODSW8jvKBbHPyNSb0rD4NCaQcJ798Pr+izvXvAu/QtwTAx8uI93
E8miYEBqBD56bqaVmwQDTP2E/QwOsS2olSgMzVpA4x3OTl8JjvudS8xlbZ5q1F1dNCQdNbZVZvxX
EPUruynhpQs4Q2RjpaGIE2T8g7DEh3vR9wW3ofhpL+V9iHzUzz748AdRYDNrrzlXfBAzoKlJBYfd
miD7vIgJYuBhBJ8Xv5fhbP8FQYt9Rft9K/vhD9hBy9htNVWFHVIwZMkMiuSkjyLmnembsqg6vNG2
wONh47kFOWJAE++ksKQTQFPOzilJQDDiYMAZybtC8UUdz/BSdHlLXY/6bc6BRA4FE5aChpma91hH
dyZ13QgG/NnSU84se5lAAO2y7pfheDklxDo6twQLL4mDdTmfkBeaK+5zbWirabzP7mBJcultijqs
qVxzujGnNOrAy6h22/21j720SSnSbAaeWn3vy/OVezGvb6O98QqBR05WgUmzQS7ftKvZ2uz/22hP
9kFnoq23tMcFC5qGr7ATlAB9Y+oIdKzpyW0O+lJ8/JeZwMRXkuWc8MAlxt/6gKcuzdaLk0rrpdYZ
WTweMq9+mtr0XXuYXbd6xS2zS+MQeeliheE2P34RUTmAaPaJqHrCoWql2oVDVV5Pw3HDsRghVVui
dF0eNpOFB0v73WpzybrEWnimevsmo5K5Ou6wM7yPojN7tPlTKBR2ZZL2nKiP7axY4LvHFDDRvJcq
zv+Zj2K8O/hT8c+wHX/szM3neLGX+AlzTSf3uBbewQwr0A8ZnmjigB7ucApIOvPbSVrzWCcKq8GR
4rdiAulgyA5Z9e5o/roJAfmdQ2wXVlCYPkpwXh5me4EV4u5MceOSmM+8vedglSj8rQesUhGFKntd
caujGi1GH9yvRRCzffm3VmLDO7Wyuz1E2OWFSDh6Ac9Dwild7ACbLid0iRFiJiCtkur+YamLXEht
RXBo5zhZ2aemkqEN6S2toBrdmBiYSaYLg9+OG9KzTpANGCqX3vWXjMNmZCrMsQlwJNjkgfnYCmLp
OTAy8q45xoMHuHGFf60EOo90b/ognWmOnN7LCzDJcrXCE/kpaExXw4EpoRf9zIfvMNbJvVdaJb8D
iK8N91Yi5bgE1kTENRmWOVp5lfa54H3tIs190/K7hLQ8SRfDPcbD6Uskehi0/z518gbq/57RnE/p
Q35Q4VeiYWgX4TiHt7/wgynvl/BnBYT7nk11kEG8Z4OdHzqNsbHEM6RNo4qumZA7+SvRtgWpu6TF
HdRXujqTvCrzQcaXKW6fqI3kKMerww4SYFfM1gYnCRVfNNBNrg4aLbHstwwNlVOOYMMD2tirw47m
5HJ2s7PF0H99M10neo+zBXvW03HlwATL0Fgbqe6FUxUnkj86V5qDyNL3Ga+SSZNil/nkPQvBhY8f
8/hDsU3LkxKiQOYq2EeYz6V2k+t7zL7XLHARTshJJ/a2W0ObVmhv11L4gZXZHIHjCisrjb+9Ioat
0R5dk55Fa2rYrKuNvbcQw6Iyv5vK/kTMnrstTzZVY8bzLyPlaVIco4rFQHh+yqS0S/+mR4pY5qQR
NgIPE3tjvcNx+N6JkllMmqc5t7Egrz1yLvJiOvuAmLky/iyJfKjZDwZjaxrolb9x/g/EnnV6FTi9
MSwULco4Gniy3Bpq9iIKwEXi2+V1YPN52Z8YMuQsQb1ymIyJKwOjqfrOKCdtf2wbiNbNW1HuqXbn
cZDPujf54m151mFe4KqGmMku0Vbasg1fLIDVvqftmvBNYBjFWZyK4ghq2Ht2rBOA54/II8xAggH+
Oz+OER7OSCfe/N6RpahLFIHYtyUG9jtAlncZHPV63XMu6EwCV7jbJgljAwTQMjp9FrWELxGX4lIX
oyVWosPo5mN2XpbLdekwQBR8UNA5LdvY9yxXke5XuuYA3XzG7rSIq3qaYE6D3ymwpJ1AJJS7POcT
r08H0HeCwaEVIXKijYbyOJeHQUUEQclFNQ/eKkhyETpqkTClR+LoMndPW1NmcsZNLU65XbMGQLca
7tzM30HxvWP3OWgl0Hvyspdfw8ow0HPvfTCcEa1JK3pG6iLAlfrcp3DCEiEkk5fobFfhL1KiBJGQ
7TMGan7g5dB721DccZTrP9qls+d7cIvobtkafSMsCCGny5fr4sLbzYysnPN3SmMtML/T7JVAxqeE
dtMBZTGHEii/zW8FlT65e1nheeJ+Wh/5rbuh0VbY/4VEn70MnUEZy+K3foyY7sR8L1v/Q9GXCL+K
Qc42ybFgA38hVeNOBoNQeXcxgbhtqGJaxGTcqqPwnk8Zsrn8uxZUX1NDZfpgWy3djcuZcpU7ozv9
iUhgqldxlEEY3o2U+AghNWWbfY+humlRSB+b4ltFoRyUxrAprcgJqlfoEZrl9qmBHiNBekQ46rOg
mQpJvQ8g4h1XD+ffS9U10RGxTlHC1CkBU94zRGfKE9RGWx+J8MiOJTW00Wcdaxifi6oeRC6YsQVl
lwRZnE4SfDNYL43PdfZiBXrSw5apTwlc+ZQRFI1WogAyvJSHsVML30ovly6guD9hy1QINfGOnJAO
ogJ1e5zUVx71jrM3NUoqkm0Zz8OsQzvA3bM+Gbv7rh6Om76ncGjCuh6rjpR0BNJnEpj/7K8rgvAM
hRyrawDutFaeCwKB7kur0I+Akow7WwynECwJzb3c6VE6YDx5fAQM1RJpytrQQvIlvBcIXqdlcNmS
0Ohf1yJnl+GbFc5HS4Y+7ydCrAZmIizlFhUKT+FEPr8ffpXIL/xr7Qrh9k1Gqs4corSbM+dXUBXc
q7GlibfAiZX75n7MGv3DW9U7yOqlFb4HBOeBVxQhwnnEopnEoeIRL7IEareUep9gKFajmXo51xCk
9/YmmSuhr00anJn9KybPKPDIadFbpHaS2XS8U6J9qTvNl6+GRY9CcpL0Kt9Sl93fR5iOfRwu9d2t
FmzPYkqRCMoz916trhbGQRdTpwJj5pd4iTeFaKWzFCK99JyPQzPWgUxooxeMhNEwDvFISiegtwhF
t8ieSfPAQsDTh+bLD/mR0ysUnBIGsQf3q4rEOhXwVbRYJbV75ihGxM6YOkZz1pPtzw505YeMQMGE
Ls8+ok+vTTFzdlAXX6tOs9mf3D5J3GRYSyUvo7ZLYJiBKe5yjpFhja7s0IDsNVKAIS1whhK3gqvF
0hAnBFTURy2JxgI2Sn62XUx3x7SGtuXO/wQIVYziAuzkn8woa8gvBeXtzSNQ71eEfgBC6XTaY0BF
hfxE5t4rC8LoPc7CZziEwnZZc6YMEEuU2eRhCyrOjG7al/MM6PCP2WrMHFCLQQ7VrYkWkV9+l6TA
/8ZXU5ByHuUKGw3jftGoiIV8uq5U+GzK0OAoC1aQJCP9oxf+HrNDi7jPuU5+ZE4SidY2Izbz5MMt
z/4UU79fXDT9h4WKAvqmSvlTs6f2oEppSjwuzzP+gS7sFTeD1DwfCGWyWBUZm0aF0SJoxtNVGk50
erLbHok2AL4CVwUcMOxoa1/DyNIIC7lYbtw8R88sEX7XAl0MRA08FgBhsNQ0MAlRp5zxRoZeQtvb
Vgixoy0LWSrh2DpUp0VGQoTGmzb4/bOBjS2IhsTO93S0tO9TrMmA+Ah0P8EcXSdw4OnlbVencCvn
5zLlXY6gRaksfRsupro20DSASmwWJIeCHH+nlyok/PFQwznDhDA75StiGFWtE61gpBegcrwuvNWZ
+bggVEAW9rrdO+sfbVf1WCpk++5MPP5rJPLBnjse1ARhEdttU+mscI+iZVl8puOIvUlQkpETxGRS
TFM9Ab8DM8lHnxbFglgFuZpg7VBnE4KZcsItZciKjYO/4N/yqrbi7gDOrw3xZqFuHbjZdmV2WqIZ
k0xqzXsFWLczfgRMHEyvGYDviI/71jYCx9Z4x8ngfEZFr3RDWOMBP6Czr50nYrlbpnzjviiCWaRB
LILHT0rG1pmWv6/eCqln7sqPX4aWb2wkil+halp4zyRxVgKZz2KgwAeDUlckCVQ1USnsTaTnJt2x
P47y1xkcrQ2/bLEVn/Ek90yltf2SESFfhGuP7yQu/E90wHNcLNK5OMFU6rDbMpZENoqJAtrHTYCR
FBVOLa79GZGEofTssNHedFIIzNeh0+xgTwF5OWs6b2TCT8K32ALjr7csjZCwY0VY6eEFKbKXTWDC
u6XciNHlYgPGXrLVUlR4PwXt6pZD+H4zktTHAsbJBVtdAvQJ8CbdyUVftXzdaRe8UFzpBhBU6RwA
gJXNZn69xr/Vo8SJyqY7jVbesxrh1HGGFIape1Lq9nTgqC3esGvaAcLYxexcxX+yvhbo8LYBHLy3
qcj1ednmN5zYXe82G54QTN+E9Qm+xoWygW5L6l2nnRV6EKfRwNQWvm5fYmnST6BDuQ6CBpJOyyBY
FYP9uDIqRR44ctZxiSiTwLCPITtG2tEW41hw0mGeI6dTOz1ZPGG1D/CCyC+6XwoYlXkpRVKtb2s6
TeSPIHhafHCXvNBEbp4XGYcyqMV+2rLkgNqtGUTAEQFXdP6sQBg/mBR5HKSr95veirX05JIk4hPr
gRveI4mRZPzQ/XVZv+UJk2Qv9SblWDxDHcRMR4uCJOFkDVg2fJgZKJ82FSyjuHE/z9QyiE3GpkEE
+p9VFOFk7WStq3Aw8v7uKQJG8Zw1h431hIpxL86ROkO/Ssp+ARW9Nx0t7xe84f1U38+S++Drj3WO
mRK7IOoLnLPUx2o6yuaINxk3vtlLspoBQErNfkX+PSm+h1LwLX5X5ZqVAgupB9ZlpFTyAyaXxbKr
idlEaLp0KzpFirNnxkZhZJ1ue8wnHv5SikZy8jlwbk0Gn7Ja5cppSJchmF415jgwNwd7kOxK1iGx
mk1qvKap1gLHClBBkemFxw9xObrzZy0KkVjqdkcBlqn/Oa/jn58Qg0CErjx8GFMzjGLvCq59q/WV
9e5fHcNLLSvco+pnGAZWioZzSlX6KvLk9PLmGwQYjmTV1Vs3g8XD7EI+EiNRIdBW5YXTpBc66WGF
LNE+gjLhE7IK2yYvvlM6v63bapPtmkc2V6Gp6WJqfW6wyG2bagQon3KxsM51ZZ/3mnCwUGcZMT2n
o36KZxNhz5w9CJX10Ow5Z1V0nMPqwv3rTWNRONAekPd5Adkw8GXbc/Q9K0fvJEfDvvPQUTwHbPfr
+/usxdhiUNlMN9KzYprBUqTFtmxO5eYMMu9826vp0VQwJS7JjbPzBlvMyGbjASwes51QKalGr+UX
ruljLDHYjf637hHtOgbOGwkEuVt2MsdZ/xTG/veNHBY3v3oAAQhqiHfAcfTZJ+t2Me3d9bEeAF3s
7TkjMpdxIAcmfrBOLCJC16T6TzLHr/4GuEA2UkBxCCA8tZur5d3pd8b4i7BrzdaLvsHExNo5bkZ8
pIOGQA6DykBgdhVenT5ZZGFsC/eoh+DYivPEPa7VyyIfmYFHGR4dd70v0yr+KHrqWQC7BqP6o8r+
9pTi+DyItWyqHUDSBEIP7B6mr5wfw2o214OLADD599BM38hZ+rxDuAVLdtR65VwipKoqbJjCkegr
yd42ZW6DfSAXu7KLMqzclq/slnZT0IwkStKxGnSnHYDJm1z9EDEYRbKihu0SATp0WxFf4DX3vnHG
I5KC4XHVExKevY6AUhBWpYGYcVAOpzyp0vpE4TrxbTDBSyXtgpVvjWOyAaz9p/konGM+ps4k4u60
tn4iOUD+WpEVl+kqTfrysi4UMHtWaKOUsYXnqIJbQZvdH2oH2syK193n3ITnO4nMCjQdPw3qKaxt
zpvt7pc96pEu4pPVHH0l4Rv3qT1f2A9SYRPhLxu1FKhr7CwSeKsjfPebIsp0YaB64NcuzHgz2Ls5
io45WaVvrFInSJQR1xpqysisu1LgdodGqVzL/DWQwx9SEguR+l9QX5jxVE1adNB9pvD+22f8fnuL
O/zUOK1zOcjdP1/xxWD2mfRiPjVW66jIepe9ACzWuapDHuuM4NrfChj6Fuyd7EOixlnynR2qAN4W
98j8cPOVcgb58Z2pNnmQehvDE/TYUdgV7x5EadfJO2+G9QcJPrjaCgr7XM6jEMPSxm2Tvp86gL1m
E/HSR93QJAEiEs/em6IMFwj6rVgaRh4XJrgRVh4mICiR2M7sMAPNSIaRBRnQF7elEDhMjqOimTXe
VVNg7Rv5iJT0wH3hOwYMiLfeY05yeWw1knpyouc6Rpv3QmyU2pGEfatcYYoIt1eUQrhCuDMBeP/E
pTVR/37i8ExPNtJhG7H9hvZdeNQJ+aK43BTiYTSY3Mzp1QeEZrt4u6pDuu2NA+n7yzqRHsntkbtE
k0oaBB7vcMZyGgjXm7uIGTldNB2KvNtBbNW2wD1Ml0lsp8zeD00BvNJBRjPVms/2gx9zjE//7Tli
2DbgX15jBR5o0CrpayecdjA+4NtWYlKwpGAbelxCNCPsyEzCXhIuFwNSG7OHrX2m+6tmRWM0q/UP
4UXidVV793roE0n97y+ZonMy/FENoA/v9PSqLDhcsu6w9VcdX54XjakrswXMBTTb6wTFA9AHkH6j
stzuFX7V0n8WVOpUfRpHoxgnNTYp52UcPAaaTXxYgO4Yx13g4juezczXYZn2YMWjkWUvGV+e6K22
NXoSzN+uWlR3kvravMjC5bRte2H6+yANDYg/y/MoMIgyRXInnIHkekzyE4sPWa3mXzWS8H/DURWq
I2XdRLN1jAhyRUVn2XyIdQFv5cs3H7CzazUb2ztOBmknx+6geanzsdUhK5nH9qpkxtPqhqeKGzkN
t56NXiKAdCqZyFUNc5Ok7vPlVcPKVu56zDP4hhY64b217wt3PGuO81eS7GcTWkSaC++DlygED/PU
dYwyySTEu9meMdJH9hm8PTvJBtKpsrB2aCtLj76HfhZzeKoI9izWfSulIRDya5MXAh3auz/jmnuT
CrHc62PGhcjCCZhz5no0ATloMidcn2W/e/uF+kzjO8Ml+L5ouw1vSj5hLzJWPocjgUL6bAsVYdzm
CPb9+GHoxKSq6Eappj7L7aqvwxAysPQYYUndHMf19qtH2r4xfMh4LCiRNK8557G4uPgGCOceD3Xo
dGIv6evgCSm1QreGaNSA0br73gnVbSJSjkilMtLG2bf9hIPGxRj4KWAOcD2Z6aspFbO877n7gecz
0AwKJTBoYfaJv1lq6HIrJNZvOPsK8ZhVv5QQPvZr+nuMgxtKrQMwptk5VhCyzazer2TVEAsL0TOP
yOmcxqRltj5EVz5/VdmibPGZ/3YSzsznmnpoc1HuiNPBVF0zQj84RsFZaomxzQcbyU7iG8j92Em0
L18d48uKjR1I7HhKW8i6eG5ml2+ibCemhCEldOKNDlNDzBSjnJWgoTg5RTBfC/pcBKkzn7cikfHk
RY+A+gtZWYDGI8YYxpYjYc2FmbJms0dl2aPlYBuAy4StJ6/cuHVMGo+28cwCaMb973ZFGPfEXNdv
Up7DVMBozeLATko6SuomQEWFr+8zDlZIQUXLwPg01/RrtjcAOCDAVj4T5u9376YBCekFt+2lWjUN
8txRC+nWbsc5wyGbdVQEp5Usxu32uwdomtiTL5EBOikqvVA/zuAQvY9bXRQhty5eUSeXsBlltqPZ
1eyW/JHE6K4ikdgCYLwBY6GLrx0XxIBPwBpu5Visr/WLGngR5BqLa/lZMaYEtiPF4gsY2i/fOsBA
ibwqFYCSoxaZHPWDuesuDNQPhKPUfbE1cv2hWzZwwKvLt59sxaL7AboRaZMFr0zXQxDUPIItcp/c
ZWvs04vU+PEYegk5DP5isSI5Hk6LRGuGld66j0Pakrxk/tMQkFSLnO+/pHMAT274Oqu4lxBVlQgG
BnWfGE7ZvhZz5Hg3Hpxw7g7KzApPW+P1mZXkseT+fArzX63o4+CqxhyVURqgxfF02/AYCJtFpoBF
NAeD1VU5kQY/KRSNpSfSCbuTivnqthekDa7Ar/Q1fSxcp0nWprNo2+reDcO2+losw8TgaIfjoqIO
3vgyNkmuWNF1Qq/iU6+ppgFiCMgh9K5+70qaFwdpPcSYUlbs9vmKsyzQ12Se1hL6Eyqtu4q0sWGM
E963WFyzMnqjFRUlfAPe/TJ0AxBgLfZsV1qH6x/77tSiOVHGcAi6m3sG6XWCxz0pbtx1WEYQcKlN
VZL35BMLZFRZ8Em6PXbLDvyk3FS3GZ3Dhtt4HzKjv8IG06hL4IUf06xJYCGgmW79fGUGaNgDI1ne
NZ1EgiACN6uZLVEMMsEbi6oKDVDqZA8SZr2g8k67oBi+Npca88pmdrkBmTwGy0wR/jicGCkG1ViB
6oDjQxhM5d5txZQoOJhop+6dRNPjd60utGDSrD58KRKOGVc0ZdEp7UmDwjNyXzqd2xgyUN3+/ta0
PNOXDdaBL47Pe4EPzGGQQenZw5sPXvneQJQbwQZ2rGbuIFtkIeegiUX5SiWg66gI3R2tCveuF3Vx
F2a/r1wRKIIP05F2WBwnh1Z4yaaoi+WcikZsdcV1MD8bKIo3sGdhyqZ0FUWmW7aP3EE382cXQUES
8TrNS8pDgLPuAIpiqJZmtVinYaN9YMCfMk9ZMg++hIUqTOaF02qRM9c20f2sk1ZYltVmecRSjTPe
+EEw2wI4v3a0NM8St4+FQPBi9ePkYPi5KREOfFr1un8Q/55Z9C2mTSsh7cjDBrQUbD7a/Qbor1XL
b6sKWW21wxNdVoMn5nXtyrlqKQL+zA2pbZsAb9YEFACWFAH6qwUWmsP5MJpzigs/5VeHA/FeGAij
QqT9hE6cddeI2w9o+inHHyKXFExEKnTq9s2RgLFHRcGW0JekFF3wjSU/ckcp0ZyCm5Ay4xtKofGU
fkLCjnJmd1f6UAgFq71Fn2QjtYNdvoJ4INCOkqjgtYVH9s4o+SlPaUPWROihiWSIJtOe/pwFSosd
acz0Wfyf9HhNPqvkyDYMEqOcOAqyS5dIMdfiBW7/3TmEDeB7MUEDSyAz1orbD6331C5FllDo1SMB
G4KqO76O77YF0XTmiaPfvZ2wasR4opBSG4SAcRouQiJ8OgNOgMrpzI2rcdYpwHRn5vLXWr5aC+8K
rs1WAjWLkUa1fqo48V0pOHJFJc5F8NN8hw4KMzVwEukPVQvwPDlAcFIC7GiVY0bNeR7vzO2EpyMv
or5Z6RDpgPHXff4rlImwk5oVrMLFHzcxsgTeWb83/MocpEq3cwE6uRgxmpAaX6tC+oQNDnI4TQro
kcsDUjQQWEkRUZJXYh1Cyx5VBDyxpqqsQ+yRhAyMofA8SagBguBrE/Vd7yTdZQi2ZPEb/fzDQ1QY
5PzqlOd14dfR7voE5NkW6SG0tEvlpYY5iylWJdOlBt7VSZ97dSsUQ8leVO5c0Gz5sT1J0pFS82un
LaCd4Hstsdw53wK/ebnY3/4fbkTT/5F7lsi6ClXh5AY03r7eX9740Blo7DpusJyPMooXUBPx9hzW
sFFc+xar1igUqu5nrE713dIzyBvqTlKv4BKTbYtSGO0ZFRgW5iFK3WfUQPiLn8jKWlyvOdp89eKE
bMOEv9gD++kyYijtSnzeaDLhyhQkvtOX+GP0WsyAx8qHvK16m7r5gAsB8Go1vXVHRL4TYFNolQFh
QsHd1T6C4txukE6XH14EgiQta72H02y6Z1rxh5MtXgm/uthOxx1RiMao5u6y3jPqjM5mYT/0JcMb
Q1T8B/hROyYQAb7AYGBGY+TsGC+yjMC5g6azUvH4va9A5uwLc+WCkqLoZIXJfSynGAGP+O5rpXl1
PpWpjntQD3F3X/qaKTWgUgYqDcpL5IS8aNTkl38NreysxQms2yXK6iAp6MYzDjTmCcpAzCBSZpJh
9+YwD/f0RDnp+tkl41CST2OGkfN2uHEM8iRvkHHK37rBe6l2Y+W3ce3ZhZ1xNyPXofihBMRCbdvO
kDiC4bQLyvXSiUfFud4MkhPd9khfS1jErcti3il93JXKqyBDrtKDHrsCpTd32vUz+NdaBBLiOgSG
pQ0pzVrtK6Z5ZdkbiyG/CchUcdPA9o8AOFMMkhERpIr0ffSqGhhtOzB8cTnjmWMX5Y5Z65aTQVL2
nKOmMp9491gBVrpbwkd5rMgHpTGOWId9dQMt8nGZZ3JWZ5UAfM2uOkfWedubj4jhXps3PrruhW9H
PimfmLGb8DCpl+S9bufGcLZXZuqKJ+PPD0PgxWwfhwszYp4YpezJeQfxc7mUD9jd1bG691FerjYs
tSlL4Xcbq2AyqExQUB2BotrbzI0OKsXiMBToHoO0pWy5sNESUEOGJp+pPj9xKDQBIKZX7r0LoDwb
2zKiM/sFE3LqB83fjZeyz6tdqQUlMv4+Iwg7KH+VbIUlwjRwp4oukSc6W4Q2TWHzAgG7z6TTfXiN
yXC3qS6oojBxADoAK4iNGxsuYWV1nfs1kBlb4rwoVXx6H0Pq27yoS0PJaDkMm1ZEOAvR+bPbrSR7
jHsKwFKtwVVqEZqDIXcyV8elsfbNLLIVv5eC1UAD5vogMHhYTdyJx5qp2sJybfbc17t+c/HbgNuk
91BRkVKMyE6+ELp9XGESu5B6ncckVdcoCYl51mM312kMgl+M1+dJoAkf1U3zIrc59eljw9X19pqG
ci+ZPyWPdSOhJEXdFcjp4GxmwzJyDo7muFmNGwZvAGk46kn9pPaA9Leq/HxPRsrKASFxvK/pNLxr
PWdgnFmFfRMLFgxA+8MnACfKOA9P1CtXbl9aBpZUDJNtNrePxHUVizAHPDnVg401g1TdN986uoeK
W4bH7eM1M4stlLrtUW4S/m8xMlP/1Gi9EpdsRkOxzBPZeXu3BjUx5Es1kVQMdA8GcOL3X7ylS0sv
pe/mVgbcK24TYiKGLbfCBhDVZl6JLiRmgRjtfVNDeO5P0mwnesGEUB9dXqF+O34NlGV/jvnlk+ko
mF5ARV7LqLtdoVwkT5C515BNSuBcKrCGZAjkg57HfX0sO9EzWSCZaYl77mMW9ewo4jRDVjI7y4bm
iNY4WDcVBgjyhTAodHTQIBwIM3t7kOn3VPUEXy6uRYUOJ6DDj0iyok1TJDC2yai7zGL0u2Tpy4HX
PTkhn/Ge+TJPoSEFKnipOIm048s5cJqFajN7+K/E9zOb3lw8//uS6cmuVsmvz6kftmLsyw/NlPCY
W57pGZzMxQCC1RaKELiHz1iBRHcKE6932oob9IIJyCbuzaH1IN8h6rZ9T5ylczv4MMeFBEGoz6XP
KYw7pnI1d7SsJikQc9cmxnzghWgo+Tke5eAgiJqOgQ6Pse9QFhgwI4GNr3+ZaRkUyJWBeJRvTwvM
DlTv9XaQc2vO+t/1SgzPWi78aLzPEcLTGw0SLp6nMl0CGKMNavdeziYSKiriaPH8cmTPeb6z4k9l
Wsxm3of50ESvaRaTmcT59NiaZewe4UeJs0s+REryENkKBDB0UhC6G0PXiI/dSq55N7ZI4PF6s4RU
J3SPJkf+wxSpFMRjI8nBIaYm2hfroHGlA3hi9aZjGr8XQsfnHupMdymf9DoHXH73yDk7BGN2G4Nm
AB31tVeC/2CCoENXcegThjJd+H5lypdCacfzmtRrOoQGF+BRDreHDISxb1Mel87Zgsf2BAbrioX6
1G8WvaZAr1EBJEfsFj+uSYh7ShYkYs1Q+sSI5aegFtA0RYga2mViUsuhjNAp1rXE7HvnSUYF6gGv
pEaW1WTYU9iiKfxlaH3d4jwHHRW3smRrD6vDEu7rhUwKvNdDxifTE2TUb/giSECRqTpvoJWljMZP
82dAobefFzGZUSNAdxi6230tDWKWcvUti6IeZ8cNpt3JuwsNfhyl+CFCQbed0kDaj3xdoIS5GFEW
l9NIE0WvxkOtMIUtsYe00ZiNF9fw8ELqU0VFGzi1X6GCjB7cok5jjNEIJB5k1Liv9hIe48hXn+jM
WLTYzbVxqeDusbpUpSxbTpEg3aHCFbXhv4fd4GcVdoVztU0EpBNeSYHbYRqJ1hz20RTt2DO3svEi
ThaJCBpOWbNb9AO+lcltN5kujUteDw7nMm1F51aslrjNsyGIujwZtjOpoLzNi6FTzX7rHkKLc8Tu
NPXyLLyHYflmPEQ9906EruGdsIkOp/TLXiKHoYvupYfRdC4MqcVjsxWM3rfmud5cBGknfLAhqRQW
cP3tFXOLMRdKQBk014e05yNBQrT6J677Ewmf9L0NoLPfsBfde3H4nw0wNTcXSjBge8FbQaSwN1rP
qIMdmKKRJJn+XPmbCOJD2EsN4mzH79IZvl6DpTFEruIzqe+DKnf2lHhnEY6UGsAV2m6bXwntZwVB
rZnmrhQhBrEult3IIYmmDZQdkwQp535nyk78L6sWSKyLaiRPpAexNXdRf//zJAgSnzy0dfdWndjR
o1w6heOvxz7d7hWAhiGe8JlpqLoGTKRTUyzbX33csFJMu39R5HZKmYL75sO4GesSTKDOj1yP12tm
PWLOMjD2wnjLbuCn1RGyFNyi1YCTeeSxQDyN2zAcC0cDdawgXVVIvG1SLlZM3oDGJD9oqDgYEjGg
4ZrXKThAmXCF9g5YXB4maK5jD+dR8ukPkNUpczzf0/rzAWxmxMiuO7phpWEZg4uxeVp27cu3R8Cu
U47AwoPRS1GTIONbPakTPaqeiUNpvb7fUb7giln4YnNBixuMdrV84DYrOv59u6u++0zK2qYZ0QC6
j+KGGEBF6NQterHJnmw6IryTqN+G9NF/JDYgH73SkotZs2XcNWdhpauGq+i9KmhLOppWqHKSTycv
4nsPjCebp2Ox0DvyVA2NBs/qaGI3xmIyISx3T9Yq1HZGohcEK0NDw9cpYT994i79Et/uRFLLe7zV
1hGV0mSu7aNTOD0HdwIiIBsEWb99t6HNa9BmIat3l+T6pAH/BgNCb4b1zLwHwwsgA8Tvqw4HXJpX
F8y5aGkiUGVG2ZeOIbcY2n6whOkZuQdZcOARD89t2QzAzwSyw0f7iiZcc5CGCSKxy3j/P3uf1s13
3KzevfmchzuUVfHmTKx2sC7QBsIh/5p6K1ASPGTljJ3HbH45oFrivdm6wqC8+ONaWb7TRhDGuicF
pVt0CtohGg4z1OznvdjQ7G8CffZjgUNJKGXKjJieKgCseDZ5vt/BXEevkV2LmkoMcu6J7lTCBpOe
cTzMBT9mVjfbHmcSzstmYEHFBDNHWskvjUNzD271+BRR2CWlZKzvxIO6FCbq+ZTZz1kuWnpMKerx
kZSBslGakuwUeb4RJ4ksAsCksEk5OxHSezPa7OxArlrCIFHyFmml6yK5lHYYGyqH3a5tKGBhGm0a
zMJPZFL6XwXAkTtNilcFIliSi9wy8axNRuYZvRYR5JQwX1blFBQJkZtDfra70p3OIECganzw3NKC
EAqNyJDAglRxhoFUorTAYd5MvgK7VCw1Oynx9FB97k25LNq6odwKnGZG7OEAwWtcUIbUo7ip/4bA
fcHybnKTXrcVPBvbN8IfOhJJM+cAIPhPaPkVMk9tCvrPpYiVp6dmDMYUmAix/pP+VVkIK5WRwXKW
SCgISu29pQitfzJCoToMoJ8qDgZROR30gKugLRyprhApT2mvSmJl0oporzPaFhRUn2OB6P0uEWKg
GDqZolBjITJ0oau6dwmczDp0HEFkEfdxH2KxihjNcC5Njqg17jGsIB86crrZrFq4CkrOGLoNVxJw
54D6FfFDWayJf78aNyV8hRX4CqPyM1Ksrg3+oTysnj5GmDzsTB9Mo95DBJpdSLmc+2Pq31IJrz2m
3RI4AQAT78j3ya6zXubNcIHkGpU/PKdxLhQgJsWqpFsVh7LKfRA6JYSlDNi7tAwtQhDaw8CTKJeo
S3Z6WXYH1KVS5cck4j3b/UdpOz3GTps8SwQkhHZZ5wiIKHpUqEO/PzEhFEzEngjBAVWnUAAXNuF6
8mHWTF7H87wrZE9xCIaESE3nPu5evQxPoa9BTmRMuDQpsBkkEUNx/3kotYkisMQpzeopq/tUAZQk
u/zjUWJI5ezwpEnHt59yCslxR+iEb+IOEYNEPDplI5NKspmqDVdbtOvbC2UDZ6o1+HijpUWyMHou
NdvtaB2d5neXQO3wMAA8U43t4J2XSyf5Fln6p3coTbrifV7EVmxn4GKLawWX9rDKVnhHF+X+qMvk
OEktQwupQcrZcHcBZgFNHEMq0FB2nybJMelaFJEwVchidpS6D55EkzBuq2n2j+0yIUxdiGGVdknA
1hEswZ9jTXDGOUP8+b2G7ppsLERC7K7oR1mw8veNa6y5YIOJx3Uiyg1caH4ph80L1ugDHiQPipdh
nFYe4wgo1VNM2HYkywa+G5kfCF4OoCuV8egK2RhtbKKH6qW15qF8ZWPKEXRcwkAgUCO3RsKJ9QB2
VkpqLhXq7g9/HDWULUPBnWLXFxzvUVNm8ARo1WGtTrClGji/4DobHKRbU6erm6p0wCglAs24eBNL
Z54Z4KPWnOY/srbVFN4EnMeUAB+idiwiufjlXOA5KZ+ugRJkAXSt29q5B7Ki44goPsFesDp6+lpC
fG7vfF28Ip4cevFrRWDMqFwnuRxtUm+VGnqTWlaa/4uWVqq7aONjXvmWpz2T0wX5fwokvPldUvKk
Z2ipf8LxHshh6BUJQPP6z3VJPUoT+FDS8b+1ljbblDL4cq9Q8BKBet0m6BTXFMu9sty5fpzfcnI6
XwNdEaKqA2mvGGzx13QQG/IS2H7p8mghyJZNgEa5CzeAov4ndYUhD/b7IIfl9ykO3Rj5oiX6gSW3
FdYYgIiKxTW9R6zE1xURBM3oUBiKV/nB7lnfMFZ5L12plKWpxGTCuCj/qc324PKhZNvm3HoEV/Br
iaqVFFvoSxatANQs1O+mthmDsVqzfslw/UDRVuQ12ThmQrBBOP7zsYRYYUe0mCYGgb0mzjvgKxAB
gCMlOZrgDRiMd0H3jvsqdx+lg0aiShehKXFK7/2uP+naX1ph2oHFSfj5uEMHaqX8Li7zDjDml3m9
Ex2leZ6gBeZFJgMPDKMzrliBDJG6YDPHxXeTkYXfr6osVF8TZfyhynUroeeJdAfcMSLtwFp2QEs9
9ZlK9jFvB0yLeEdBNhL+s5BVtBxix7ka8fzc39EoQfQVIf9pSZlcnC4+brprojdLriEErWBDFevk
66pqotl5niBTi6vinCgAIomWNLRGb8wbA5m+LBwOgIDe9b9wh20covs30rRjhWs4DkSOvJlBxjdZ
qM1Kas7iGhcLJb2ZVbXOJn+gO6gwRk+llUBFadNeoeWEGBRzMwp7/9Nq8Q4gSdvYaFpxTtwLhcbX
3jyebIS7NDDGY+PHTBlXpBh+8BtUzWTaAxpi6liZOxlSrqNJeT9PFEXq7PXIaS3z+xUnJcPis84B
3SaE7AgXl28Jf/Jun5rmAq08Qgi+FGYD9/QbfjG3oR6k5Ej03/av4JOtyDDkXyl9GcJw83YOfEVl
Q6EVgMKmZ2/MBPCstAQsC3QGGkoq/X8lK9DbFyVFYhNVwK277QzRjTeQj1PkicjwSGLHjZhhlDPd
yXmQz2M3zrSkynIribkQK7VVPUe78POvUTNQ0xWt1YGbPsKbTeACivvBW0yEfLWvMZu9Vfx4nGkh
Np+ZmtzSTwFwPyb10hmGHej17LM9AYW/JnUI6CXwAZKx1dkGZFzJJ8Q1tbBm2cd5efD/aaXY4lNa
UhVO70X89BFcxkIgH7IsSi1USy9aAIMdmEv1B748X0Oas/hFWTkLsoPF/U74tRMcTBx0RGWBmaYx
Sow4OXZO2Oy4z4u3tPf/ceLhnB3R+xfF33xi4fAI9rSjYIcU2qZMc+AzeJZ9lc/VtjZgzjFfC5bj
qzMSOOeZBF10jtQMnprhhF77DlNRm6jc4LxZ2GXBf8Xf/Kfluw/KxfKxwSLrRoqyho86/Eo0FfBS
C2PErE1GcpcIxI+uB4TjVes74iS41a1/ZjgEHUrBu5x03FIOxpflQo0558gNyXGeo8Bkav6tdWuB
y4MFB3xa2rqfbiO2wsCr0ZP14xo05y+AWP9zAT1CfWrHcgvq6fI9KHYET96nvAxnoY0oCyXiC/C0
EUih5GeFTEHlN7f6KwrfqFw+lX4K36G7Jkso/oXRnt9dzcyIN/0VDKwj4XGnP2gyunYAeZMf8MX4
XW1QWPfrI69mGgWlAPOmAsQG+rN7TNb4MbST6MVhy2z6XtJHsjKezEN0zlFCYYWQeJSFRIAylw4T
wmLcSQ5G5HYFjXVuyKiCS098/l8nNRZSEiIg7bqDACaM5aSs1ryoCfiKCTK6cIenmVqzdGAfDwmK
GH9E2xhx8rNIJyNXhOskbkqq27uSe/jF9VOcbOoOb380ziAs19Wc3dlTeQxzKCvCrpqzxjudycUA
nZmzqaEuT5NQS5vv4nOte+QKbIzrc0E4IPnPueXo3+8e6MqjlmvfZfQ/IQHcCHG+a5OFFP2LQl1d
nQJJqqdlS4ovVFcgybRKbllu7R0GLzWiU+XEiBtC6Hpi25KvzBLmZhrEgz0XzJbh1zSklinwVGTY
eXZfV0m6TCvOzkMSRaODATJ1wq8YVKjObUK4iGm0fIynmQjhEKP0qp6a8rXGArjpQegHFqyA42hS
6RPwIPCEU3rxwJXJ+6JYgfCJji/WsEaQAUEGnPmpR+xKYHFnPOyocfVTBpiUOXIFFF8vhcVYR0IP
WptOrQ4pM0F5lgzAgVkYv0xrCqp7d32VjdHgf8VRPiBqOrzrv3D5AQEarS1tOtoEfvnt/DkMSU9d
gAckTkmownyg+2LoCwH590ILIcQWUP9u6Q3YTr94vtzX1kwdaKypiEFL2o2xpFCzXLmUjuVUNYRN
Ld2CNxBSa2b04aggqWQyar8NF2jTtXVxKuwdC4YsBrVGL8H4YK7x+m6Qr0V/ySAaamQo/9hdcMcK
uCqwh2G6524txrqhikfKkbIVAgHNf1IXI6Fsx277d0RTJgHIXo36g+aGQ95Cai6iqcmE4MuRPcKF
kN/eZhKEDLV7zssx0oDodq6pUJ5LuPrfdGfsyaVuCA80psJDRcWUCCKXsZtHEtd/TopnRTtY7Xjm
Ukg0ity6O8uYqHfXui9bWDjWLq2RSjKerFCoGWDQE1J8Eko9KVgGPoNgDXEYJi4rUL5HwwtTNqBO
c4vynrFl+Uui5wp7Rf/hwPXjfwikqUDLzdPlGvxzKxH8Yoy9T+YzU1AbT80e3eMLKdu7MDFi0vXV
MI7JQ6jOZI/eSFr4CBAlW3vhTPFr6Wi3DBuSjFZAB1pUeSOFAy2laHUlGVBo4uqN5xv9ITiaKyPP
jEYIA9g+UA0Uky6h2bg46oCol3f5KfdOfGUZLCfFZ+rxWp0/AAOZDGPR5ogcRDuQfkQ7FitRF+rq
hUeTZs8/D2MrwEKSGSoLp2LCTh+Q8sXcYCVPjyWBRHeSR8oQ9YyTlaO8m9vzQocjMjVDIGH1g2aF
yldX0MvXNC+AC2wPBGUqRe4g/T2LN/Q09VVmVaovFAhIhEDwRM1wmkQ1pGeECpKYc0t/TdS+nn15
us3uMT2oBfoEsbJvnGw+KUmsbO64tSLkFl0U8xooxe4dg4zXOKexwNrmXE0uT7URR5sFkvhfNKFo
NFqsKcTGNRG15IBHC7Ju2CqZcXvaihLG6yVbJL73a8SHUEwAP7FEcnVRnMVlJqauosH6n6Gjv1OO
PCVsKIN4KLg12lcu6YsamcA18nmy9//LLFOSIK0folCGbjKRrXPv2Lyh8znN3eBsx9mxU66MMTFL
C9LnHSSPgSeu9NJIpcyn73/Bp6uvHAa80P/FRwkZ7iU8jiTkZdKaU63nyTc2BJwuUuXSJpbVb+Or
iHSX9xhREjQ06hpQHsAlFvonjCzfiK9utRMB3fTzDhSXBSmfEDyc/SjBGQ+zGFVM62vfD6ww3Z0T
GHj8EneuBOBaW99Wxm/rJiy3DhDlaubrh1OemkZO+LPae8gfJjIvrzPFsVgsYdNCjPKg8z/FJCXB
ldGRVmGH0IYKWPKniR+3s2pz4slgVHedEtTPjl2pyh+LOYonUF+44mJ5sRZfeZqRC27/8ZcUnKhb
uFEnoFM8tXzYFZg+ZHkVhjqO5ifeUPWIhF5F0uz8ECJjepzF58sKXZaafI9YxyYwL71mZyJrEPDg
5ZsLw1mFU4if8yeD+quFI6GbyOT0R0j3ezI2D8EE5F35WsNu7alTzsYQhmrcDe5GDqd8wOfsIjBM
19iWFm1dlG6WFFMSpJsIIkowj80U/YsS/l2DRKWY/n8gs1QTGj1fldZ2Etec09h+u+IFRPn9ZRI0
kF923qpyTJr04GLlC/LR2d6Eo8QqZWZOERkEzu2mwKCCntr1AS09zn+PBYtBhFpzX/R1OL9Htu1x
WPvkR9isFirV1S3oK9gctZZT07Pe6R9GNPlnQ6g9RP7X0wL1XPgDrpDTXIpmW0efsoEKyrGy3nVg
+iVIFSfpXkyIDY9Ktl1RGRh1VAzuRmuFr34XUCYRno9NOpaU06GqqcyTsMT3UXHE82huIHFhegxJ
QI5E50/DkIHuR2JejgXgZhYVnVltW2my8LyZHiRMROxJ+Dx+PmuT3Qt07W8rrPeOuIjAoA60iF/B
UrlcBJyfmMyQZ0yZPZSqNlHKoe37PYaphh/YojVRaH2wuiRvC9SSg2n1lgJZLIlMFKey8eX4eBhq
a9Xs3Sbz7lCHwfesE61GWUcoOo5pOWgkWl3hFntSSarLgyB72tSlnugvk3ifFBqjGHm1HiQd+80l
8uuBG2I2fPhqetvq+NySHQlVzE45dQSGFMHsokfXH7YOn6v/rf0nIXQe+oegLKE3tBAc2YrsVqGy
khzR6/wGnMu1yV9J98/C6o9hSqf+k2HDykftziLZVBKfIxL/yZiDMEyoD9b5S+eHxqfnVx5spLhw
V2G98irSk6XKmP6xiac7lcmaHB14qkkTPddNZYuTceYZdv4nzNiwANdIaQQpakcx1TVcW9xv/8Xb
xIMW2Qx/mFMNYpzwJTgrGHeIc+nzObQBcqKPYoUKGY4BP4Tb6GAujpc7GRAMZ1srfvbqF/4XM7al
aBsO1Opq4JID5uIrBx/BQ5i0M9FC/MMDvPVqSorv91q1Q6l63iGj+2ICN86sBaSbEk13uxVM6QCJ
lbieunfD3bZYI5tOHr5KuhbbLoG5WeN9kbKDtt0nmXGibUC4lAHaKJHxSv/ghOJ9U37v1Cri9A8g
88vm+jRlr+BXl2dFVDHymy1bSMhxE5qkFw4GohWRLgszfWItP8Ybz4AnM+6NM8ILUmjuDmJaFOrK
lU68n7b0f14eaK0jh2ffXCMIpJtL/kTM5HqQlQzF6NVvkTc7bBEb1aSI2Urso1feL77BDmLOQIOz
pOV7HMeKirSV8Y9VbNEBornuBrRHMpowJ4aNGNhl9nztA+9ZbQZF7r0RQaZ95bXEUs1AVemwW2Bk
DPALroVIhb+YhPbKTzA4ekwkTfazQF3s+xv6wGgcj/z2ChCZivCuPvELVtDZ8QA06prFGrtyu1w5
Q+Tfw0NtxVhekmCB5QOfpddwpLejVCRaTSD8SPecGaOahlAeoKI60IolN3f5K9H4m04dNpcBi6+o
jl1p2M+I7txEjNXrrXcQUQJntyRzbGMyoDMcKwatlqCOpViv80/Vnqz0KLeD2I+Ma2cWKswioPaD
6YWQR+AWJA6Ty3zSazsRP+pdGgn1gro8WCTIq6/2lfDKs7ZLmBcvWa1Cldyo7WkxuaV6If/EKO6l
62ywUnmFME8SZsSxB4VVJzhAbW/LFInO8Cri9esHoVVi61wU22uY9mhvtUbLwmgoXq8+xaDhBmRt
+Xo4DybL3G27Cr0wQwSSf9TOP2ugIynfxQ9cblKGtJHp++c32+UlepK80gX0MGhHp/JELwUpClFQ
gPYlF5vMY1Plr2AYh3y/++Hz5gFaQWSTENXkEGtIUj01m5RN42XOwQvREscdBiEDr5Z3gGbVTbZw
Sm17NnZUpBLFQAXDTDcDsqYd/HoRxcwYApti5mGH+jn7VRoRUFRbCv7Awkj9/8IfAjoYm80mhlkM
IAiLRKtdSSHMUOkVTdIeJMGcoELB3V5dIUJzDtxNqILFfXasOyXikQV+uZ2moAOjB8sUYVtFp87u
pip+ecGiNAl6JMIKgeIEuDXcMhLhSDiKQjv3PZDKeUv12l7FUd10HyXy5LIAjpkqjDeyPVWA852F
KL4lMYnUvW61J7yi+Sm72HBqtuZp8hokIKcWvCao6S9zrEI1X8OyGNX2bRBXP34tt6gr3M1g4tdx
QWJWj0HytCJPkA1KKiccpDS3phirssheTswu/4Pd22ynMF/bYoTmcxf3rebfe/Vx95Y1GJZ2zB4c
Gf4el4n0NKAphnp8OcBwQcyQnhobjCcp8OE4f0DOP+0ry2PFnk1aXSm0Kcd9qWk5jhiUC/T2jFrp
CMMNltPtfAbkmsL6FynsGriFiVMqig3E45sseGpz2VEKMZABZ7j2+b4x3dwwDUVXke4CnkyaCG9U
oYkCd9ZuKFX5wy3meSqll/+RbyzdZFouC+jf+rxMJmZ23sQSjnUlIJfVRbA0EX03iOtXnzFuZLXy
M7ds7l2eGjayHB/Be8TMtW9Ngc33WADObSFlu9AU9Bvxm689bflt4kabm/Ze6+i99brpuOaRGmfQ
1/YZurGxSrXbuY95vPJwOAEQqGDos/e1ur0mHsQvovb1tfMvvMSeVbTMU7r7B0p7G3v1SFULE0jN
TapYrkqejwut64NcyGFduqrT0jK+mkgK+aITTzNc2Z86/glbXb3LQ0lnCyPNVyvBz8xrW+yiQ9fc
kxN/FJgJFH5Re3vxOdiNCuQ6PlWyvJH551qoCjXHZsd5lH1IM3/xWMGiRmSDxBLjhdNpT2z2fACW
zMZJRU/neQclg0gTOOJn5XVuZnGbAHWnju9X9tpV2lQK/Mkn1XCdM0YHulCd6UXfxQyTxmphEaFR
rXHYDjlMwOORCo8wsNmv2u/liuICYskvJyf2OhFa2dLN56+6CHO39LXUgoY3mqvSzZgd1zBAPEHV
KLU3/yflUBDjdYiUYcFWosSqTOywjy3jekVkT6pmPqcxXK+79EkjvH2vfS4FiAKo8LXko2Wgpo//
H93LcKH2aSWrdEHg/y/vfhBoDiq3WkspjqaGq1uKrOAMbzfH9089PLeTdUuLzrstwnTmlawXEU1t
xz8pya0EXkxdadHzeqMaqjoGL4Fh0x+KC5MethAlKKvqFxPAEiaDlCisafNzhdYMQksTmS2lMIGj
41GFX+Y7eiUYPS+Ymoi9cqMx1ef1YCWr8k2t98PAPS/r67xuLKAi2n3ny8sw95dXniqEtMAhNyEb
ndIgK0LQnN28xLS/6HyM/3/w0eaz+iSCv5l7aB1mDrDvHxyyCb/FhipbmWYJZGRciaUgimUSRXTy
+IK5BiyBJ1vfBLfy6IwLr35gq++WAH2FgbP5pLXSDVmizC+ZjHHsxkX5BIIE4j484Z/GjIxKZSKC
fnp6HVpBsVH5pPxyz6bikG2r+BMsLAggpMaGA4UGRmfpWiQp9IOeU+n4AaheB7+Sw9hd+RxiNELL
FsyywwFGXtkkyWazSCwf9HUAVyGxPrScexOrR7Jisxb+8wSKiyMd9XGAi1mV0853Qe4/9J8R2846
uoEvjJho27WYMF7L1M20KwRhZ2E9ED5fGqcJduXvmGmuVQm6/Qor10WjQAH34SGsosUODs1MhdCZ
Tc7nGDIXTq1I4PUOk74mnpCdnS9f69TE3k65mZeQYpWKqIxk5zMq0EGs9k6Cn1bEWCvWPaP546+F
VWXhmXq4Kz0aHHlBlG7xRYx1i8S+MTk/bl3KlR6DLmZQCyyXODLK2gi4yg1te+sGj/rl0rG81cuX
BJDJGzfMoNW3HQoA0Pz5USLFlzubyge1Lmp8DZBvmUcT7ig0XQ6W1LJXwBhn6xXoGi6KO+rBWBR6
KyHoWqi+Mx1WxI97Pmzl+MdLtevfi074GtDYn6lzuGjbhqanjQ6pGKiib02HVqkrYLnrZv9Uva2z
1yvpUeRDFojgq+Oq6xDw7/Z1879eD5pak8qMuqxw/0BAJkFxudmLQxbKGnczcV2Gq4rjhiLFxJPq
+m3qTpzAz6gFJEUV1/kgYVJ57s0CVBR6mIC2G6+Jfi0Tj1YCi7jYmCrupAHVVwGYDu4P7uRH2UTN
t/DmMhEVwcS3IXkrAP+LU4onQytaNYpMyj/Cp++8vsulDZn96aO+YomZ71/UnxZimIdnfE7mpocc
P+bt14r9HbzR2abyLGcIRhdxLfPnsL2DBPPI+zLnEzS9ytZr7g9+AjiWF0j7r8hwyFIz3YFr7jwC
85kFw9n8zEpWS36nNmEwGuP9F5SSywTeEt7YZggLhLax8UZw3+yaIbRLh6Al3rKiQcyNP+PxqpaX
58YMgn/+cB8IcvI25FsHtJBTZSxsIDHadZ8alHys5UEel2Yunr4ROmCSD5ridMR8KeMsGrOYylye
p/McRKKLCTbf+GRhn8G5t7KXQUIakugrfxtoXDOqU0koLFMSPqbQnsAv9uNiOzhnaHS1i7ivj13k
VMT6E3lEpzuhcTmgY5lFdXiZ6XRzHVVIQmfWKZ2dqd9BW73HRZin/KybEOsJD0+5Oe/U5XqZbHH2
DHT7njR8l7JjR3yReaH63bwO0bl5dL5/2eMW8NwhWuuPgBd5VujJ/kki17SuaZk68jTzFwdBkh36
LcG34iQRoWRFl2KSPVC4MYhxmcmlCUWSWb+UvUeswaa7Rok+A1VpfGqIdqAqkDc7ze/4udZBSFTs
2/645PpnGRxbJb1RmUPIQP0dzVO8rsA+SXd418yBdGfHT2D9gyOqBYMPd9uvBvOl1OTVNf+pz+9H
bIcYy8bhLp4LskuE+E2csHJLqYjYrDatw2WpPYO1hznO5m6CMIPNFohLPOJG7zZ7Mhv/KTxOBxWF
c+D8fplKHrqptL77Q8+xpPr7+tYEcaUxIGOoJmUJjrVGNUzSto6wlL50gxWWQf1MsnURgw3ypNLY
CefTn8EYxsU8W2Z6Ckv2N40K6JebPkJAcgE5Mj2cpkYFtwGbkH6qqkqzK0HHYXt0sJsFNFOwuJt4
8AZfUTtmHc9jez1BrQYMwHuydW8vNjEuiRYUbVkPLBYYS8ArU3oCgVRCDxW0AzIfZryjHSlL6JIL
nsPMJ3x9R4RI4im7VwWMuKEOhF3Q6hx5IbLupbC677wuxS612l7tZXYF+9yHGMPp6243X9jyj0Hy
ix7Jmx5lT5XsFI1XkQ6d2AynzrhpLl1p+2WPZ0rKocnevFd+43CBBsODNzDImNvoIshofb9crOX/
J2XJBE0LkR6GFKHZRm2Sll1X8MCECNFrKwtIJSP+p2eNUJJwzCLtexoV8rjfvrMD/D3c+XevbV/n
O6L31x6FNRUXRBc6JaYS9N/Ps7xe74JDkRp7A3ppoZFP9vtVcnJlQcjcYMGWbZ19/zpGHCYZLKtq
3l1sIy2kUmf4+YrFswJNs6qKk5Ho5yzEW2JRFwUFhxOQ9Uu46/9OvgtNrdNShoWlGEs/zK4gA7ce
k5bzeK0JFzpOrrAYr+UMgOsX3RwfcYKVVxZaWAv/vR2fM0R6bCwj+lLVFmEoTgJMoFG4SeSXKk22
2lvBZAmW6fj6i/3VxhD2A89QLUJ2nh0bHerHXdq7n0oZKttKtJmprIKucqnDyu8KPngu4TRUIES0
7EafWBoRuUM5G18yHnO1h/CodGMXNiPjVm7hM1kkG4hKSFGHsX6JencFR1F2igKx2YySS55KxLHA
Q3RPvuR5wOzA4ky7kx2NDv1g836CX+qqmdRuw7f2ybdjC4+QJ3Nm6ITyUVe/pbUu/61zggeH0AzF
z3gZjmV33evgqvs4+96kFK546YHFwq/cXqEz/9W6m7nc8L+maBqUUyNJAzKgXkqSnqsIVvZPq+QA
C7NmnSL9z43eketAegp6DAmgu8ezEDCZ2rjRfpvUyngw2jn+K1E+1G5GN4RusCMiE1XjrcAMv4e5
VH5bJCiKuqrpKlu/fQ8yYM/UZyMCwhQQSpr/uAfq4JQ3ZEpzxpuoUW6xEDa4ctfMnAgwQSUfDhhj
Ugerwy5YPE5dkrFLEKAWbWcDDUmW07y4m7Dmw4e/tingS9pwN/0vnzz/YsMRelb8PD51F+Y/wp59
QEDl45yxJ78NzySkBAB9wTNXmr0Pvv6oMhDaAY4zUSjbmTqoFyp0/CagT6sGLBmX+4n+qtZ4bWHO
ru6Z+7Gpj1KtfMEIaWOOUp5YYk1ZTbIfXbTlkjv2FBGh+rGV1OX5ZAeE6XlRmiSWcsvK8P3J5qmh
PXRZY7tBN8y30GCWPYgGpzdi6H4jvl9MIevzDdSZ5Bq7E3E7FO1FxRk+Mn147MwwLhuy+HGwXHPF
haTaJE3f7p7q+XyBi5i7BVJsiQngGWFTIuP5ACrvxbSLa+2hWjL2kDdu9vZ74/VC5jISRaW8F+4/
n0i4Eo7TzIlHy0+A8hOLDB6eFdEyqck4r1WpwNKUZeFk6rdR08Oe7O+JLEij99/e42VAvdzk7JWD
vSURSOUWHB6SeWXbooz3ODqVjzpONziswOA4opPLWPfyXBHtYyGouDQxZGp1kWRstm6AW5D5k6vi
nD+b6zY3vgBgI3zTVYWGiUsFpZv6jmTzCIfHGTh0lYnTB2MaSByujpDrNv+iY0lvD/pXwu+VxiJa
YYH8IiuBSuWveTIlhCR+VfFnV7VPr4H/RP72rn55Up3jVyqhZUQ6/6XZbcoiK78DPM4+ce2YkwGV
YFsocvwDNrtyKPdpSK4EwV3iY4WqzylRLDl4Hm90BaldnmY/HM0cSdsjgDZwhMASTdDHfmtjzo06
sMVAU8Efuf8EmXcnS2me8RSYPxGgKidwRm3OzubBozvObRiqDDMwVCkH2pKd87cVY5/PDhi+BDXT
Yivo79bQnzhCas0oCEey5kC8qzMjQCa+msOzFPncUyj8tgxVrKN3qx/p6o3epKwmJdpNfThNxmXI
vZiFZfqoIqAzYrF3RIVZ27JFa9uSmal9OaOgGJqaNC0yyTR+Ygdy60y3XQGyqRnCBtaFqiMzIhKq
1/8DYrDzv0TYMQGKxSd15Xwm7m2hnof/5UKuEAJBN61Ksq7XP8bi5Trr+rZIb4Q5ivg3CmywNwMA
BOcWAgYzZ3v5CtWHBNglMwodOq3OdTPLuAFGxOxMpmHu+D13b0zcYDVH0gaH8SFbroQPSEotDb6s
w38fk2JoKjgQc/rqlH3GXIUm9a29RtwtnQm30Ri7NF+f8w07bOwgmTHrBqxyZyHvH3NzAMMr178n
HUXn12aW916HOTVbgXlsU9trgF2GUfNRJ/JS21eU/5LfjEiKkq/H/WQp9+JSepn4sM+BCDv/Mmga
b2GlR8ZMDtc9i9iBY8u2aO2khR5+JgG+K826+BPuPRZJFwmVNxx0qr/JXVblI3g1kkQRNvpMaoY+
gpEWQz+VKWC4afsT/xeDCI2sw2LL0sU4I0oJYS8e9o8ZOJTgJ6zT+dsAfOpciGZUsZPGFdvHUQ/G
cGUa1JQYXZSSLyaxmCOpCjOnklQA6C1t/4QOorhTb0MKPm+AoDI7duDZMjOG3xKRBImPdFwHZTux
AyQBwta23+4DAdO7kc+pQSRMK3paOQOz8bPeATbQeY+5ClBnFhzH7zEtsstS8Fga/98NiVMofKWr
iPXr3xlqs23dYQXpuJuhTg8Y6KriEv+uiRuCkfBVdaWUpUoYDnHCPejpTyU1PqSKeyoN6oqpxoA/
YXQfIKODc6XMmTWy5/gisyJU10mN8WsxwnGTh3PbXWVDjk24w7NwIrLuEakD/DGRrbtFqsJVwjrs
SRI//hEJal6QmYkD3rDLojLfvuZjLMrCHL+iT1LiwqkHvh4poVUFDleb043eSKh6copgU+IlBlVK
PRDOfUNJxSOsxEdMB9ZGyENPQkfD0tRJ5ydezzOMIZpFPtqU+wx35FxhGfk3qrEu0M0T/27V5W4X
IBk9+nSYD7CpJX9gHYYrGG04xaD6VI6waGHWkk1IAkWtXmcpq4HBjeHFh6M3g70ftmel1kAqHUPW
e85PcTZ6Y/JnDcIfEUxItrtltA9zlLZuSHSWRyNLu/yetmrE0YF/idU/slvk+TkLwo8zRgt+XBOV
gTygL4T4YPcd46JymQrh+MDmwVwZO0Fq0nhK5PnpM6z6N9CWGjtck2Uol19kCgIKoYGLNvqwV6+G
My7AxQiSAyuK8CvLZ8pSqmnZq1uEUKMdEvSS1kif6iqus+nqzlwFuv1h1uyh43Z9g12dnTrvIjTw
yciuUgX6y2wzb9yIifoL9UkazdELxCOl0cr2egen4NP7SJR3/wv9a1zIX+nEkWhlE/alipA/3qNA
9zp7qBzFvAxS0SVluwslTkLxfqSCcE9xgXYqSzmq96kCkeF7qsjlQp4efdg2DrYnesCWg6bk9zur
wARpd3hhuNmTtJRJaw4YVZBkxeJhPKchYUYYpw3t47ZFi+SKWOivlJNgqn/dtiB95JtMU4uSCfIp
Av4jm5dlcmlX6qDo/bZc+kTnTsoY1GlSiZWlHyqdztIMTRyMW3rQz6JyTR44GwtV0J5hRGh/Z2L2
apFQNEG3Vl0U70niSSWtBSUm3b3Zp4OTYgDpzT2569cFpWed6duCwJWFueS3+m+vVjxp4R0fmD7e
LdcjbGIbgnmaro7x+VTTF+LLxez4gBiadXH5nT9j447CDNBl9x2XSkr5cqJKV56xjTQH8Qfxby/6
49dqaKC5uF9BGhr1q624/gTRCBOqaw3L+nJp3ow1Iv9LSkfkQoSCivpgUClGitJCChu2yjbLri2x
2KicYhTVbC1nNvHFXFTo1s06FFH+lteYWdavrOPdqZMbgQERcf9NBMmT17EbQL/x7yMYGoj4ON5F
EyNbnM14R481fC+ZBj9xy28OBa46ZyF4z7d3Ari/6ab+nHHdg3oFWWRdRCIo2KJum4V7vIVXfGpW
rxPYic3G1qXGHBIWZQI8zZX4PTgU3n3ZBjjI9ySFyUc6KmbFG0Wb/eXk89PGH8nrALqE0fnWx+SH
gtFMVE4ILInVIhVWwmadYsIahYIQlOiHAx6/nZIlpNr2u6Sk6po//xZAd7iRKOm2f5Ob+UpGFot2
HPsgqOCnnjDK23jmePbHgrnBhMuGN2JeGjM9yi5L1YbmrXsnLWmqrhlbzsKo7cCkoORwcIwYGT5z
1+J8xqpcNJlEIbZElhto+k37Ce3UYRlb1y4nNFAooq935DYxyAE68dltKe4DsXehw2O72Yb4KcAz
iaFwUdARDgAyOaUJGct+Rjfspt8UxGsaAyrzOzX2/f75l7wr76uilYfUAkivQ6bSxkZ5Zw6zf0we
Bj2F2HnV+x+u0vheALkx+tXJYsWBKW2jzcXQN0vN9xovP7Nezli8qfjP5clbccCCQJ/RcuILIYxU
lPLiuuv+TkJRjQ/RUmm2lFYgajjcEx86eyQZRHYggqAW8MohLSuxlIXj5jugNuiRuxL9p/7Ee+F0
gT3U7nHldmmUiHRNENjCW52CnZlPHtAAphK8eDIg0VJNSLiuwZrbxf+jf1yoUTNoZ6kk7yrFzGZU
xxmZaop6ah+JXYzidRZhf4ZpKicTzU17LTsMwip6Av1Z+gWp31kJAY+PBExBYBMkVyzjkseMReHd
dcds6ceDlyAZeNpcAjstvv2T8xwJ2bUJ2bT4jshqQYy5flFPttahj3+tgNSNEsK9N4XBOpyo+VxU
9yrKp8uwB1OEMVN40znoTajkeJ6mM3n2wKdtgfgGKnbnbujOY4K8dmnsVxCUzTc6lNN6/1rsqHmU
Pych66ZGBOvv2ZCttCgfAkAk46wZSYtpGmiUqzkZRkRIUUmnSvaqdoOo6QibwWm9HJtl0nGvji4o
mvOwSkigvXxcFIU5ShzvvFhS32PSmYZBwpIj65EmBvHJMUsqU+4g6/dG1Eif5H1c7qTAcr/XgehB
HWQidD4L4rxm33yo+txU9wsd2dAcavv4MuKIjfrSjPmbpiyImiXGUABXRIWRGIaPpEYjGf4vGdue
PxPdozfsONj7YCMNsMtyBlMuNUDVtKoRijTOfqoCFEe4nYD/JVrkEGU4n08BhbdSlM+WXbUqtIhf
X5rbvmja8dpIeZNyLN/DdqQbt3oWAekxLefSsqpwmS6ARWo99mQ9mumt9885951wev7Xs1+p+pKr
CDMU8Z9Hfen+psuQVjwcAD9ZwfVGcVncc8XXzCnL65eKifGxRI6e7ItdmGaIDSBOIEE7iIxG/hVF
Nx3Xd7SA63DvtTxRIfeP6AKUlH5lJX3G/cIUGlRrHSIN3US/I+Hv7rNuMEryNls6wbnVQb0zfk53
+A7qB8vIxmHtOnvB2bEMYQMzmhxiKiQWhtoC63HXegwvO3H4f+Pn+2Kt5wtUxnMCnoSHG/ckC6at
HifTKDpzwb2mHM8JYQkM7bLsP9QYhlHrY/5oguJFcTahnf25dS7zofO8SD8Djh7E/X06dvYP7Ovs
am21mqWZ4brjG1rQQFZfaRTg9GlBI1tUtLfZccRxlVYN/C+HNK6rbJB+dDJbA0JRUe3kZO+p0xKY
7YJOmas76sO7q/dDAnxje1O8/rEjNZBahHzGzAWqi1dxBjnl/5SUgSfGZL4ZA59vhB+Abcu8Y1wG
MqwmHRPxa1NfNP66+V9r00ysUFnOUwIZQ/8KO6RmV67zUHmVfbbfFh0XzwIiUr/XIUkhPwzpfta9
1IJECifEATHCWjXMAR5E7Y1bhYG7oq8CcrUXF/NEVrV/Ub54vyDFWriBwYcgBiJjCtaWfvxGVD6H
Z9X/LXpaLJGWltqH3CkqZu3QVH+Qa3StU9duC4WMPlllIN7Lcdadlq9nIko+HakuWRUDPlC2ygw8
0vKlen1Bf+rgNz1vhNcFslGrwyOAAu+q2IKNRa7ePvpQd3JI4XD6J3dkiTuQ43HJ+6KNEjZDKlFP
T2Ar7vifWxh42MEp1TcZb0iHTIwsAF5s3RMPABAonQNXql9/2r/IlHgi8MO1aKeUs8hRfjupf/6y
l3j9nlxFWTgMfLpW/2l1LM+RvM1UCHyLnT4r9sOipPmqF0faJK73y04K52sd1ZuLae71CVzWukGd
WaUmzIEbb35+S3JsM68O+14o1SeztAYRSUkR+3eJjoQ31gD6trI6qkXUI0gRIFpF3qOdGpKH9f8o
NVXNwALRhJwpLKobXBCyMKOqUuJ5PkgjWbo41AMF9NnIFjxBbg+2JCYI860iTLtOvmPEaeRUmYWh
o4R/NKKZq4OHQjZg8silrEBknX0uMGGwAVNnPUczumDP58qujPHxfh1Cjcgl2Y6K3ivA4b4+ufj3
NgKgugHJxfw3W4xqOvSX05QfJcB+ueOgYsUJRutK8w+USkQiJc6v+Ur3eieqsqNWqypZJqU/EZkX
bBuG2oqogwPQu6cGBs54xetcx//boX3iGUHFRDGk1/+KA5TU13NVCxtny7wv/7qBXYopolzkX+Rm
2qGMlIHanxnT9O3DjV4lrV8A7mlUjDaB8QPMZkFaDo87vwPYt8PanvQLCV3EM5hEqMb4GQqc0lFW
o15eED1nr5bbKWzk95Xh2XqYH2f2WTmgUG2XPqOCoLT3MU7J+kJBsmhLdqjDYF3kbhg/tWjEY49X
L/YfyindrV2uRYcr6woEHN7/bRFaeNtpXCyM/Y0PLhf2aqGbPq2/BD/IqrukJs38t4PIgi2F/3Ej
fnvyPbGg06Hwpz1ihGHQJq+ZZqwNGPqWa55+xXwWmWvAvPbTjxNSpmnqnHf6kx3JtYhAG2WAasxJ
Ow0bKHiVmpeszhsheNljitdhjev1rXIH1CSweABwrlY+WH7RweBbjClyTgecOhOekblKNTaD6bjq
5oMSv9QB8Uj82Ga3j3YvB9diDZaiZWC4az+vtRNDeWA1jGdNuMuMXo/zgXwnSE+zCOiuLyVhEBCb
zt32jUz5No1XOodQP9e6hNd1B1o36Uwj1k2xpTwUUmWEULfTM3L4yA6TXuyxZJ3AHWeg8krbEqgT
/k2sruSwRgEanoHm57tdQYXpQGnguPbq9Gt/UWXfqTfwuzVFlLPBAU2B6eR7Yl3C0sEY/oLizNCK
A+sF8TqnEUNOwCNV58CU/cPGETNp+0bctVIOxVTGws09si12Et4iz0pT2Zgq9mwLjTLPGB8xBYa4
xBsQtWH7A9J8fhqj/lK/yp5mCfrb0IJSOUCr3h29pt5XhynxJt1Hv0l28hQOdyeXOeYWZ4JyWAzW
pzHUcGZ4geKqBfam1oJ++jDAJisLP5c/WAi2b3+HbEJuBZBbIIp+rO/InUMYm+cn49jAU3j8RAHO
KDMB76OcL/3AFns6RASe/ovE13klOLWQv2jEiSmnkqVNw+yc/iJk3UKDbVKSzTDKcGYb3UvOVG/s
sjR2NGXvXGrgtKi4KAzyiAHt8CAuoyf3hoFQYwI1iFIRMU3LoqWP2cEsMJMioKNqYZkWTT7aGws2
Yfp4kaJIbFPHUzVlU2fS1+FeMm4Ep30Haf8QijZoRzmm3xN/3Nw7jbXBqrgFdbgIiU03je6GYts9
xFGthqVIoyYcNUIml1iacLRBx0Vg3axO6yGw5nlkbbb44PXzZeJRZRH0sjE943+YxFq35w9MEoWd
/TQWpNPD9uGIJdl441LjKCA3hC+ZmIlyVQEEvht0FoZ0bKvGRULe06F8F/xGgZIwi4jMq54Y82U3
jmyboET2cDhZ3v6XrYHyAF2B0WI8fSw/lwIE4604q3ahgd29z5bfCAhNDxwXSJJKCtOJpFTu71Yr
yclF9VeIfPhftOXXKyPP927FxMn3lyNnzpWnff/3hY1HYDqMEeemOkvNwgTQ5xexhsXsVgVM3AJv
Z2T3O1MevpVdUE7GwkcEPRsd9cvxNuEcQ9SQ6gQ4QYsqgMsxmVkxmCEh6Rfm1m4O3HQafjVrg4m/
rtWGCTsvys+tJrvZ17wQLejBsw9HvDyDkygdt6ukeFwhyhzKcB87UfUhepsyMHfvHvFjwVjta56W
KrJLqUYDiPLk3BJIf9k89JQcB/Wyxj7QTTS4/ym647jb3bZcFpsR8ZTAfsZ3IWocD87cNESo96RR
u8mgjY/JcWqX7NWlraNVtUvDIiFeU6B83+RT/w+a9JGarGazV04rvoLids+/32OoHLgLjNTXNt5d
ncuqEnSqn4c7Gs1aLQffnYleAhcniDR3lQhfKOmnuDctCgcjArDgVKbX3cMZy2VMa8FRY0SYEa4q
1hioYfizrKufpv45Egc7FivydyWQsyiwEPg1vmc7LWXUcqPULM1TIgnYbopgXAAHp2No9B9J81ar
PwhAJe9UHyOKrWqHenThk9E6juoDs3iVHNwoopN95xAdsDr9qddSaxvGTlEdRxoDTb/GARgkcaNO
wmB+kU6vnKYQOqX7so+iLMtI6n3+8ZowH11PyDJAJhBsjHwCAEfnkpi7+IoQYw+riei4iVELb8KF
KtOYeBxOUocDIl7/+OoK/TOIi6Nqqgzliytc/aeX4APAHsrn5Svk30jSsJE0KlKmDXRObehXay32
CQB6i7ji/22Pcnc0SLqq1GUDG9pDTISf3Wi6HfIciRHQ676IPNZr+jv6kAA/wGGJie3/YNkBYBfw
UdlHclNFbktf89vuJXanL7Xkjltqt4zjOcCdRc35soGlGBzq7PGCzivCAQviBPBM0cZu7RaO99r9
yyvXYwfFhfgREcb2afnHBnAVEKCSLCBAdw+zwofVxDhJuiQWY8sgEehUnZM/hZpIKArOhXYz9GZ9
v9Hk0/Sd8Q6nQBtn8E9UT2qmYLwwEcFBC+UEdrAgpfPbVN1bH627SVzdyftJgiBQ1B6zJ2lYsjCS
AFT/ND+6JWfgVpoOMMuTy5dmcivzxQkLN9Lp68kLqmC3h0N8TZuznyd9hROylTK1FuYE45QGNhel
8Z8P9iG/qtR6xTBgnNuTSupsJ3LyoQqVXMzS0owd03wsP9KMwWhhKkdDEwLZqGYX9L36nIo9WS+t
5IdqB28Hnpn8ppUgJlyrOqvWMAeFwMqtxuv+afztDQpvYv+/fSBAJAPunKqJBpOi0Skd6G1dVlIb
ef7Uy61l2KXnYV8i3D+uYNs5qMW1XnquCbsBfr4Bk5XJJ/cbYdplPF5K/mevZNccxj0raeAyfWEM
GlGyMaSIzy8nMa1LTrPkHFW9rIQOsqPuSke9C/MDtMDqf+9b1n+9Wo7FqnXmQXL8Bjf8cFgewsmq
mvpkJLMDHXdAxMdvzbmHkyvIJeTDpGrp303dPBBagh4mFwlMbBTxNCZhaVPbri6kFKEWb14sY8tN
+KehCO/2nXN589cdqaeC8viUQ0xDZ4KWlXYAjkEEYuIYyfBpXe7BcOx74b8wCc4h4/StEpEof/ww
NrRhm2WmtkPtVF9uTHYdrkxd+gO0U8qxWZgvyfBGucdf4u3anIiTbfZM8l40+7otufqjHbiMpIFZ
zew1aPCyo4QD0Lt+hUqLP8VdD6LQb1CpU9ViQbLFGkhBW+bGY/JayfVZRn/hvzTXnyw7S3UMHPVP
zV42TGxIOmBG+IF1nwkVDAnWD3WRWitWbvoxWcdzul8U5uM18WbXx53tu1V7qPk22QVcggGPh63G
0v2GwBRtjzixeojzAK22AGTeKUcgPHaUGrb0RR8VVKD/p9xpyTiGNTFfi03aNYvr6MBZPLBsl/6z
tHPws5hR3NsLMsE0f/QaqlnMqKiqPc4SKDNjvjDbAxRTkPRQhbFgdLfZBFj949CKPnqiZkhwHeoo
KKEJkvHuaqDuSwHDMxDGw8SuouixyvXK9+1Z5dDMfhmCxQnopCR2c1SR7b+ekXl3izwUBgPsucOl
Y3D0Ne6kXTBWPyPQDuyTwREkTKBJFWdVhzaYiD8yfoxp1C5nQqqRlXGBiQ7iLryZYlQLedxMM70a
xVsgcJxEGlfXG8WNS7X6aSoNud7I77H2Otm6o064nc7gf8TC1lTZwRgSM6yKP6Ryu7XUO88tV9+V
jytYIOMP+kFDdIWUAM/kMYSfLClR9JrGpObnBuRySOrQDgaQtSeZ2TFyJm+0fZk2Rm8H4UUOlzW1
ghaAzJ5/3pk2q3UufuZZf0Jo0/y9nsGnCl/fle03qSlXSYUSeQaVsPNBwcFeKWUpvy8AGd+EZxWW
OuSHXaiFChNu3BUb7TXYJqLrnl1vYTrl2Ckwt853turECZspk1UNcifMn7qBgADSb7oe/2KtqANT
YeLiyQ0ENCCF3HVTmn074rAUqc9z+dMVvTAbO1LWP9R0Ddb7j2+v23QJSq1L5GCX/4DUukGo6W9N
3GMNmq1E/y53ZnIawr8E5WJXKH1Ms4KY/pwym4ftA5Iht2u4GD0T6qsx8WHRuhgNbhEZjHdp3Iad
bfz73N5KFaECmXtqqSGaLkrT5mt7fPkR82uaRmMljlHafvhYc7EgcfiQoOJp0yE+bEvs365woKD/
C0bUeKtFi0sFGAbuqr7sTeiteqJPXsrDi72j8X06YkzPoRXthLBElfzrttP+ep+ClKpY2dF0rOfm
6W1Ts+JYyP+m+F3cKqtstf8l+wa2yEhSSPbcg/mTabVGLbxN4fQG+mHvjZzWiJH4Em1BBtnLLmI6
C5G/h1t8rHvLvTLIyFOrhbE5zsn+m7yYH9Ir4ifPpV8EdCX6W9iJXNI5PYxRBy9I4jdY3aJsJf5M
Mm8HSGuc02Cirv0YnOsp9VVdq2O+plDciz4jAprzGKxbG2yDlmuk0Y/ZQBfKCJdlGc7UefY8oW93
gJn/xPV7wMvS1cSHQ375SxoigWX/LQRGPOBAo8fVjebjaVPEzkETrVZxksgvMxQTxccZlUcep1Oy
/x8MqBvaQXiVC4HZpVzCqqharkHW/1U7uqAOs6QjY9Jf65jL8R5lRlat3rZALDp6dS2GOqcBv7Lm
SCSLWkmz4ywHVyLlsR/kZ80yXrCuqGPpQSYMkU21bGia1eqha8DsgjV8rfiRHmTkyCgEaSL2sbBU
zalUqzfefM7B85lylBm7c6DZ1kC6BDUJ3mJgl4sbOWwx99F4EAIAl8DL0K+xy/yHlE2o+SFFlWTh
9qLhi22UzSrxMPLeRB8n6Lkyx5IE46PVHsgdjUT1wqtY8BoDR1Scfd7Dp+Hswt+IvWQQcF2nViqe
/BeeZEE07GDZ7o3Yji+SqfAoH6qb49sQXR1cVgTl4I1u1diZrytkmrRPyGOHnxeC0p56JORNQhcB
v5Uk7DJTVqAoyB4+iPvnwd5vjqiqGWJLWwNQou1bwW50lmE5rXh/Rmm5C5pjiBtv1NvHIFmhHO8z
6uMLkcJ8JViurhHSXv8xmw/cZji4fsw7iPmUo9Fpkb2Y6A7K3q68QARuyBKXgrYFFxZGEddTcmuy
gChHdchNx06JLQzwUUuWaFfs5wbhMl0t6e5z8lYKMGdrdfmkfvrSgdQGsUCEUbYK0a6JguXGKLZv
269/ABTpKVtzPH/CCIDtRSdGuOG/7c9RQVybpSXJXB79RkcH5PQKxoFK36WnUPO0yflRG6YBeCJu
yB+BCcAwH91qnQVX55v5m2Pdfawy6P2l30voNDMgvTq68/a8iR3g7oDkeuYCIE96s0cByvsqJ5F6
GoGBt/4YlR29ReCdKqC7JVDUOvDWosW7Go5QjhbchFtkIET3rNMep5gAFLiB8Pqcpn8M7/Fx2c/o
WT30OPV1464YVzpDQhB+nEnX7ajRqHWj9LOcaCpz7dAfV+gL1YJpIhgK2wW4Bt/zV7oiHnjsnVuL
E1I4WE3MK+V0haJY6cJGR7pItIRJMZpBGmAxZN54awZtDINcG2uCt7vY3GmM+rBIZIkdqbEtya+E
cRsBHok076wqS0RBXfwCT/Vxv+cNDzhsAfJdY5uLIpFIfllJKeCWUhi2SLyhJNZwmj0dviHXGTwT
LaLIC5dbhBnwmNgqFFkWtM9ySQ/77sN3VgdG44h8ki7fgFgvUQ7iWTJ66l2zrT8gIZDNUBgjKmwa
d4UQ7I7G8EKUP0W9Epbp6PNq8vdBs3xJRP+sgW7hGDfpMuouIg91ZQFRQjnD+12XnWwPuB0LPcfi
y72UESRlBe2Zm3SqPHpG0Wn94JtxzlUQ7WE9qnfzCxLsGHZQqRiG8YTQTLf+XqYdnegKZW5FHn0r
LlcK6QtR7VVZ0eTDrzMNFxT8SeXUOB5C2Fl9BqdyRA4uAfBTXjoaPs5MU4fQtWQU6HRjPG4GlCov
aIoE2I5x5BdQk1pcCGnGBy8CqvlYFBsXpuZXg+HQdPu/HXs0945q9V8uLi8zouTNuGO8J8EvpQv5
ttivJnend/Dc7JKneTPJrTBsd1sbVD47gWORDG61q01gKZAMV3hkG0PDgsHjm45e2yk8qtR8frPt
BTfV6XRzhHUQjGY/jrYT4cXcJCqasRvJDau/EBJ34ujXm+Ry+1yqg7GYpI1r64kW+GdaezYL8HZ2
MaAtKMZlQrbMxxN40QVqAzPiE6aecLkzowsjQcQ1JPjJ6sxzPMixQyuDX1lR4jr+f7ON2BsrsupJ
Tl7AFKCnwoYvuPLZ1RCU/s7tBWG4VPAnMU9RgCXfBrT7O+kI+D68Dh8AF4eDf4ZvkgtCHMkI6emn
F0zUbuF4pqmJI/U5vnDGmcweE4Q5oTMUtKheEJoCAw4BGLgiA7kfFbMM1rkeHD9NqpLIcmIjjfzP
dPdj1RLIaOVpti2vL6VOmW3/y2UOf8nLzyLSJPT5Lg8viVvGit5meGqNnbC5GhD8A+znJaDWl8kQ
IkZ5dGxbKnDgbgfs9EWH4W9bo029KgsQqdlaM4uaX39XIH3Q0eaVqT7BqPp7TiTib7vq3lf/0DZ9
4H0Ulgl0JQCRA9Zo3VX2APneJJoQceXakG+7VPdwQ8noG+h2OfuSYhAYib8VuEmitzKoWUOdkanT
drWsPLfWW9MetvdGQycX8B1wpm9AJtQG8+ZsTvVDIh+HjoM20DWTjA2EL09hQ2Rx+RKFVEKTaC79
OJPgQZ6pUAW8xD3NCWixwUo0h4z8HEnKsIBROuuhzfffIH9BAvIIaOXPmLgMRg6xd/SsNa8Jz2J5
T89EVazbK4qL1ZP+tTrt7mg4+3l5fSEUlkMC1hXNx4MMUnXXon8n1O6ibIK7jhSKlVJ0No8l++mK
mYfK09xUr+CFUkOYVJ5PNVcGyxINbzL/FqIHf1m2ZP/JlyZliqoAUwDh7D1QlUJoraO68lOO7yCn
gy7b3nJxZj68TOu8WT+m9bTMnFpuVzm7BdQs4HkkzhwD63cjOzbpVzmPPDNAqnnsw/87GioEvbgE
jHyBnNUZcuibWbILzrpj2RTFsgxaQ/FNqDCW2Xpyn9TmXhR2jWa8AUyNyG7d7Xpefw7+FVb+4Rs5
80jbSGA9/M4fStQFkqPjObi326W5purOF8mY8KqUOUwVJos9XDhJ/nvtsIVKFUMC0vbK5bVP/1Ky
HF047QziUddObS0mTPmPQgQyKmdTaeTWosVfWw1aRHZVXOJ9aYGdAxW9fXtDahkKg69t9djEyrzw
WysZp9AVdSfRqvLcOIhXA85WtiMpqvasWpuPgq0HGijwBqr3Zax3OxSWQcFCzvcr1odpkzYfuesk
qA8bFFzLAxTkCR7owLaQY34GEBIVrEpbOHU6XAxSGLXE1Bg1IH20u2V2OT2hVDte3WTpma9hPuc5
rkEQD/zrwD1SKm4PoBw43BSZVmu8UYlBoq1DKbv+4HTTwc6RhezT8F7Q1pD34Bd4GCO+ScnbLqJ7
ql33V0dFoVNZ+kF8egFmhuMR3MjzQrGRdXKD3OT3OhcWkJSnckzatAVM5S/xHhbSGNZIy8Z6RSBR
sA7iHLovVfJ0a/CGfyw/7YicIUBWJAGjOtPZbnGv/IHz8Dmy1zr/H9AcunJVuc9sfYc3CrUS3ADn
Qwipv6dM0WQ4BBzxzSP0W22HDPSsWdpBaBi8XUUcFjCKOn99hlVdPpthVPKtAJjPMhTODMB0Ud42
lNmbd/OQtFDpINdBMbYBPpEWwWWRiBeX1Sq8s4A6IsKa45ScZmflIhYNbmTKxGAMGzuCfM4QKLyu
pEFLeAmhleifh9uxsJDDKVJhsS5MTDeXH7T1E/Aerf1ap4OzXT4rr9pz3Mrav1sB0XfsuZVjFTHF
lfle1Fwih4gqlxnF1n4fOb+EHPFmKAtxbfxaGR3xQs1ARmK49cBOOe+SD+TX8bEGb89DbhRnUMM6
3v3q+8u5t5IM2bI93ZVwcjuOxKnAo/hBwCQVaPTGr5HPjR7FXAEdZZHvkQlOc9sGIX5WP9fdMvnW
d5uzlk+c5MGH8MDoxVGQmdEUop6rFaaR91drklIXrpTOU13HNJftMepRrtn65sn1x9CAgfWBTco/
XvymdAH9xgc61crA6uFlRVMaOa1jSR1IqHtpUqByIRECVgHgP6SsNneq576rGKKFUkQBqSndCxVE
KvEwybsY/ljcV52TT0JsxsjCTvAg2lGSWmaCBvIMSgkzjTJp+8RfJWrG9xgjfK/AzEV2ENOKHg/U
wDC1tcQCFvHinchzpmwqg51PhLSPN3UX5KQ5Op2lqEvNouRs97Q3CSnE/7jUrx8cWF7H+DeQOf4I
rV92Db6dybgYpFX8PsAcA4VVqp9Hv3pFVGSoIq/qVEO8Z8ISO00bvC+F5gfQwp/TQwAGnptYRcRV
uFl4ZPmIHBybXYq+//otrsLFRGtdzQI+kiiSDRfuuBKWVV2+tOie+jS7s7ICJINs0hMGLYqCJKHj
er8I6LD0bwGhBfHXvDEoFyvnStSG4VoA6l3JzxA+OjWi9esiDUYaqJYafxZU64xNeGiUgqDUIdwO
fTITtwN6apnZZRChBi3jx5ZjJZlqvnbEfmIYztzoo43r4oKfo7BBpfkgk9JgpbCWfZh9HzIhNjLG
4Lk0m3duxuyp4M47upVkemN69I0wIdpfiiobRRyj1TiSRA3UOQe92B6qQ90hmKuOqzpwWqO6PJoA
aK4Mb9XlUXOjYGm57g9ch8ck3x2M15ByNE/Sq/SJyfRj6LtTXvDVaMkiS/wohmlMO4PpWB9sqnzk
0tPslihEEinrjVKUFCf4/bqBqgv9tmPDsGfTdlKm1YIw1xRmld8RKjRA5JqMm0EyRXcdH8ykC1Vk
xICfMat/mZQczl40GT60ymDmbIHquGpSGT3A2um9aOcpSH9d5nCw5fQopKl8WPQ6apETHhLaExO5
06NWVSJsdtZtwfdQGOe0yW5BYpfI/ntFH4zQZjUyUWOgI7dz9TuaLapSrYai837SM6EIAMnuEokr
y44JQIhzewUqrVqEArbA2sMYDpDwui4CQimoNxuS3pF2TZxIopW8t5bAX4hqWYgDLUEEY8n4tFE4
OVQKtefL2Cfc5tbe8DF/s4XTvpr1pinvMG/VqTw1nLG/Gp+7laG1yv0IQRx7wFuATZj2Qd9iErT4
TdtmKTijdkeDGTJA8+Y1GaHgc+5DeLdytWXN2XkiTbJMgADH1seRMUFgIkoy6YE062h6/nCJWyhZ
fBY+eKb0l2FbkWH/kx9LPmn8SntJWdl0d2d3xP0CggEerB408Bv/lbhIaRTTtPBL6QDhFJWNxBt3
kzEpdHAbh5sdLJtaLVPX6LuYDKUIkHJneqSUpJb7YDI2I6mMfSTBUEKKShM9cAZHFN34UYzOSJ9a
a7vphA0lpMDCztTMHmunzx2KqaIhfiaMW8SeC3R5tNoH+wEH/Ut+kdiz5sPV0gqXVA5hHSCe+8M/
2+KVtjNURXj67IDCjRhxhKsUCXvwy3tpW+M5u8EjEleIOgME84gHo2SCUyJeRXnKauKBLLtVcl81
yDsRyDAeSfkChtBBNm0R/mhRSD/WXO4NnutNvU39hNOQzTFV1fZx6V8pgg2SFqI3fGGqoQHzNxwW
aNY9bbvWKPSYlli8kYlFhXfSkVxOKibMmTPybmCkSdbeGx4paCY3wFqXVyMyyT0Nn90Eq0IRCwz9
Lir8YYTIcXhCbjRkAm1uJraOGd9aLFNX7ZtpQ2UyGLZEPNE9eqSWUHwXGqrT6KLxNPo0khWeHN2s
i9nwfPSmjxyXn/7OmMzyrkKMI9QmvrsFCW/BRLjnu6pOcHTH5XwTY2lwSLhUPtMdm/TetnBTesYD
gdulYan5eu4cSmrNAj//GRcDOdJdJ2fR3rxLh8J5CFZBNaoGxXus1h8XYYp/+B8iBZR1xMyWMZO4
OyXUXWbmyLfagKMyHBxAno4EhLytmSZek5g3tQYr5hLtrUBjNbj48h5xoQMi91Hq6pi5iIyLEfLF
alxicL5tKW04g/ZO17MnxuOp0gh7/XMso47Ncy6E2ameiZ8CnbGvSpTtSgnLdJ64EOZ/smqjL9Ll
I9HRpokvECPWLnM2qcahFh2NQta33iRS9hlvso1SmSryRE2VHeOSNGe/JU5CqrwbPzR1dhsmZvlo
wwX4uxWbYXgNCKYmWF9SOdtqACamaWWIkt+8Mifar1mt5oDtw/tsH0EIxK5gUBdVP8MCff3Zcp11
y8rUIX8gmWBIzt1hOhdUuOPjSAaoR1dFcYAXPAPXkdniacioigQecfhiKfbpIi+10lwYnkprCMBO
jSyhVxpAAnIi58KcOF9DC8jxxxQP9UMGQTu0HeSAiX8iRpXVztOCd3/WwgZyC8YcAJrbbYeuW81y
2sGnyR2WjmVdM3rEvvWe+JZngCUv/qEIVtZOzw9oV6+hwM1dalmuYN2R0Rbs0Nv4Eiry+nq+cX2a
15CUjicmKG/f18tKFWv2f7WLLf/RZt9E6dJfR79x4WmFV3g0zB5qez/bjzHS6INZ60sMaR2Jciv9
Bpyv9/8tYjnNQHV64aL0WONxgx9fR979cngwMjd7gEiXaYISw6Vc6N5Chb1JhJLymTVvRcHAgN9n
baqsvx5IJmWNxtJLRGLcqjTuxqqEOvJGQ0rnS5jFWZoX0+g6CAZ3LoecxB+IZnNAOIpbXZ2ITgbk
W8ABYN7jUC94UH+qJHXbQor5sFGpSKecQloovmiTszs3034apU20iW966EvQvdvODRrzSoI7iq47
5FyMmcL7uv7YUYsPdogFABRHnzvPzkDGEj+d6V0PNk/YWzQu2DxuJ4Va9gEFnME+S5NxjMMuM715
AzoxhD74WvN/ioT0aJWFXMKprbqid7Rr8a8NeV1UKrniwj20glOEmPscnuCQmcTPdXG6otAR4Z/M
G1QV0TuHuqFFfVEF1/D3TqU4hFGetSfAzzx6FeAXnAKdUhEC6eqLaZlYe7K2Oc/sPOvQOkG9/qOP
vS9xwyDyiB+fDVItK7wkq5t5F7ZQrnf1dWdSqLfl+XZow9pasZEcvrb/2Avus4YawHlqadt/EJ2+
0nuwn4fcebKkm0Gibrj/mX0lTKLdCWJzn3YyBH1l6ql5c9130q8ezEqRkZ8E0sIpWVpWXT1jY6MO
Z1vGBhtIBO2jciEULdjSVAg+NLAo7dVYcIzt6L10KWu42dvBe4+pLgasvlzV5VZxit9WCQCd8PCd
FTBlrAAbks59w3sJT3ELIPqQQ5SMZ+7BFs6KUygzzZxt/OE4DkCFFdLltG7sFsoyg426jJeR1dNe
AFN9jek8RmF1IHr+fRgtSpPpctSDW2y5lpN5c5uscNJrbkZt34RDGo3k9uqKoFsiIxiwF9Y71mvO
3wYfIjVZF6ae8Ez8OfDG3TkK7rupCsHBdNSQRJ758DLfbzALpusOa2Ofsks5wyDyY86xuJ1W1TGg
ffXZz5t/aqF91HmX/isDCrdEPhKgVPIGQeTawmDTO6PfkL9L6r95uBfQud4l7j9C0E9VKggEQlEX
KJ1XIOhQ/TvjawX6zFrLcehUAjd6YNKyMH5HzT7E59jO8h4ipPdYrfKCBGPsdUMZ/Q05YfKdqvQg
D8Lyz+Z2obDaTdGmTwg6xcB7UlisUQymkMM6C3QcQuXUuja9I7w7gcllcn3ftc+nV6cnv0m/773U
qA3Sv9do8YYLzGbGp3F0NbRQvMzjh7WO3A7NkdY0O+EQTSDnhCcDjdp29mrZlyK+Ywo5Nddi1xwV
VSkGiSay/fZ7Lvmp2WLpQZno2QivufHdutj8FeP5ii7JclQcadQj2e8ImJNn+sq4NtsL61dlPf2i
BtyiCcrOmDQlbKGndziP29X1mhxJpjJ7f5TwapHvW1pao8LDCf0S1ozoDAfjBSpjzWok/a8XHpPb
1rfZ/XKCIPdq7kxA1cthtdaozNCL6FrgmFZ11C0kE66P/PSn64nxF/I8oqyHUgoBoDah9LVMzTU2
+XHr3Qk4GaaJPbLoUzqkzX1uKgdugQOVcXM7WrWXu2tGFZJfnMaXEsnKwLaQlO5VryRVdSsjO50e
hroR9oHeZvxz1mdBdfiGsZmiDNACFg5bRm4rFZ4ONDutEcPYPosMyDfTpjfmx7voW9jA3loXWAQd
/4PTqMCpOL4E2nCI8BKB4/yhW6Yi40f9jcR6BIXwvtNBCUKi8PRBNH5jt0WaHNEo+2FeyZ6F3ntx
cNeNLxzVTZnsPOQ2lKUJtGsrBsHeW+z1yDAWm9EniqIWywh6wHKq3T7/nv7eTXlZlrbRyzmXNjHp
JWxzYeIACfYnA2T1YzhSccIyzQ9UAHwym6L+uI9uY53HLxO0/epBwizR0JlwlXgpZtkvqm1tjDvo
YQ9NbENvOCPOzxZpZKBsvJ9uR3JhyxiDLgEvfFP3S+T3buUWPWG6QxzAggoUxoWALuQW3lWmSxfH
3vhoiSvM6NHKsJX5eJu/Tvoe1gZOgI1MkXko5NOPzopXO7Lj+H+6L20nHnUiXsKG++MC6cyqkPc6
I6ZPeqqKYpcdHtSxT6xjlmyAyVKl1/1enVja/KyW2BY+wR+HiWU9xZ4h5emjqsGOMGu/BvqyHjfE
3/sy4hkzEn+3V6yDPzVN9tMUk0Z2Rzd1xcSqdVtM3lZWBFlDOfpig0RMFUNDC+g8GIN/z+njWZBe
PqMNh1HSaWsNUt639mjYLJqRxDo0eGxv0S9VaYY4VTL7cnqLGYbBC57YlcdbLRPaVjHXdu4N0Uvb
7ujzpPeOkZB8ITG46zEZ6HrYPtGsGXpog+RBcpY9XCbG1xti02LAhgp4kgoUxMfQ7W3tII0aO5F/
PVRs5hgL5Jhqe0LMkZ5ISNCs+Mus9rvOQLeVjPy53Gj7SDHo3zE/ilwomkQ961nkdoBG+niHNCTk
uy0hM/PzWMN3DiY3B4BdT8GiX9SRX8y6tHOYzeb9ctJiWo3DJ9JgEYgpr3ZF76xOt+9LDT1Dzrdu
K0gx99h6PexPrkkJHNDFLgJm0rcuBeAee2EgH+K8dV5MVoIPcFTPb3Fu6/9/QoTlkU5ATOh5M3Mf
sKlbdbl0hjT/Ip3opB/x2P4Ri9aaAGvgHyHZvzfNSbMXm/QODaXE9luQaa/KtCFL81Y6Xs5PSUI3
G/FqpZFsP/piWHEX1B0ziyvFO74jeMyVF+nm3+Je/Vdd9zAZlRlrvpuwTLyVRzHKba6JIXEjwErJ
V/drwfnNTAlfznMSJFi7rYpYVkSYL+Jb+eSNFs+uoN/GnhDE0cvTFAHmj/pm9si8p1Noyroc9Ckl
23TBsij2ARk4VvFJMX5zd1E6HMGVgtc5PAAHHyZ+lFjucQbg1KBwlwCuZCNwA+gAI50NuTURux5Z
IgjG0uJhJnGpDeG49N5ix6QteYhDBo3avJBIyCZzCm1I2OknNH6GcQMYdmTRJwKSJTMNsg3J0uan
7qGLAmlxkhMsV8R01ggYVvMu1EgHmsbRFk5heTW2g5Y/Syd5wcxs/ff2kTmmIqJ251q9yGsKXu1C
ryjWkKUyPp+du0cssZlw2xaq6KVCaN6wWWO+j47Mox6YcN2eUlHLN4ausozGJoHmPYnDcZAwM6TK
no55eB3YU55rbe9710ntyUkwtN1DK5vn9MvRtPBp2XQkE3iOtZ3qeMB28J145OOAg9KVSclvqw2u
YduD1LreNsRZNf9rKrnLRPEi5SZ9fAlf3vJBMV+MbsTHoyKGtDR63wJsBpjQpU2oInssxRfKJXOZ
PFIIkkzItsBtdBVUvfF04p0jzLCk1O1pcUrg9stkHGERMRIFTqpqoPwDj3nde6jPj0zkkH3EtpGp
dUVTQJ0XDQVAkuQ/XBKxiyB+HrePfhl3h5ZbkaNQL2MQhUk1hYA02/ld/43qs2eSbbZXmc1GrWZF
x4Z8T2+7lafTakE2nefMessyFZ1WUYiXebXPN1W99Lxks556/QoG5Md2plS36hGBxzIJSSwgveMo
zKvkz4Wh8q3Zh7dPSy9kp5J1DGyT8M0fh6JJFirHS9HvnVJDAct7yNOvTKZlBsN4jTd4okqGYDI6
pLdJxln5xmvlfrOl//zwXBLFK3EvIMcAFC7VuS4LonqqIw+ym6rj+47kQPAIVcx9s+pV5SigAvri
gYRQ77i2L21Rkw7FwybnfnrnO6FGaEJCO8lFlyBTZHvM1Hv1sLElWDmudphE4e8x8aIZvz0r3omb
QMaBVIVvIOJ3PNxM2vRblyUBNZm274xwzSaLUJwBeEfTfqNNyP4opMpqeNJxgHItoCfJWZcey18Y
0xKm59xRh+NbP3kVJH2KmLsW4fPiNBeX8vACCy//TQ6uZKR9ewo+DmbtwMBXvrvDfw59NIF51ClQ
DXzubIJQyYjVcMfTgG3OMOfPZOmdObxxIukJ14/3ptF+ekYe2JCNyQc31CPtD63LV0nwTTg7gVvS
RmktRJqhUPDHnZNTuRjhy9O+GbOiUs1UcbWrH7Qvna4fhgGWU3d7Rqpy5sXgcoicRWVbTHrv9p4u
Tk9zlrfAVCsN98izlIcyW4yyCtcjIEH54MhvZ7lPA26cS2PWdGqKNNOb0LJOeLPdLTygIEGJSFT0
X0k9XoOQWUSqgRxI1fwfJFfAwVDP0h7Bv9tULEIkwuyQMFQD69cQb679ElW91UCdsxunIhCFiiqa
lU4K4DvuD9KX9yiLw5fZzcM21WWmK0DKop5TFGNZ3R9H6RmmXXq67FuG/yj2skdePeNjJW31NlFL
Lp7/wEdF1fh9My9Xg89x0zwFJl1pJ4JPNzXIZ86FImae2pmy269/QgqpCKEQhaWJZ/f3Dx4uhZHw
kgNBG/y53JKStSQCq0h5FNS/FIUTmXX5EnzMg+oD78zFC+ZhCg7AO0e3ovrmcyHkSoNR9ja3qurP
JdBIQqz94JOHbAQ15ld5IUxIBMPN3d67L70ILtEv352H5HbVcTJWlLn3JtEG92DbJtN3EiydAJaN
fHNh5Aw7iG746gPutC0I6Xpez+8B6a945b1oDxrHOwWFrPKEwUUHV8Q1SQJdddkz0CrH9xRvQs0t
ry+SK6vaVkkS0XXOLpIjnB1bdR7I2cqqimEE2jwhWt+JyCq0Q4FXCKWAKlxCW4V7K2a1G7gApANe
hjAKw5VaBYLgOr7kWAjpWRghMe0g2qTXubqK9WJwKFYSM1BY48QLxcidwi5UEu8UBEOJELwqKDmZ
N4UxLh7Z5Qf5ShYXDIrm7Ln18sXwY6n9rkV2jYbk27Sf1OPlpOZmXPmpIhUUGDdPrYVy3bgo2KMf
rwTTHaSgB398tXMXdjFpjzchEYOBuSJ5PtF4DC3Ks09uXONA9wIRgY89BCu1O00FNF0Wxnf4tz3T
RHpzmOJN4BynLar1A/4a9BSYemGrK6Q7gPnGpXEND9jJ/iFEBucXpVnZP7WhzyRVH+39JGFYFiut
KuGmgvSBRA1+N7YKPRjC54Qopi2wVm81eAbhJsUvMx1DpVCtYD2ekhJaYw/84Jl0SYy3HOw/oDHg
qZV+vfGH7zbfc7NFxFmZMw7JoE79z21DuZ4piTvKZYRMYiInnp5BVzeepn6qDGYpkGpVPxLaoenn
FY/X/bVLcCQ8tv6WAnHxdwu0SgzTDZbAzNZr7TRTNdJ9zGB8jHmous6vqdx7N2LUylli+29sx7mQ
oMa72URpI5muoODFu/90K0j8nDkO0A9U+g8qknhv4uAunAFCxxSMSDbt+5nylEghWyNv6f6jQvxc
bK7fbNVglTeaZNtOfgKnae3JP5IjLZDIvA9CrBiWknnlR7k0Vpjopl8VAPb8ZoT7oHVEUl8KRCqx
uxzCir7RFx2fLAX290/O5/Og2qiKk5d4cXckZKsVS/5dYVD5McHKdb+OTddnpUdQ4/Euyk+LCPWW
/3Rqf3ZLqPKvf/hFrdNaHx6K9uZMKrGfSCsNLr29SJpr+EOvPVrgVRtThiiqkTCj4Xv1lzht5MXH
fdW5909JqmhccSebTCFqJfi9Dah98GzBUQQdEwLdYY6R3YjBUEjrc+CYdyvRlCSG4A5P4VBlfXo/
i3ga5D9Rmao9YVDV7JJKXb7AXJoEZjdq4/p/0ZyVSlx30WU4hIG7ufPiVknRx3lzMlovGxHEORG6
2E5O06YlzVnP02FFctz2/gajTzptyr0HkVmPcwi0x07kD/YnFoOqCiHwpmVmzt83DlVjk1MY6fml
cz+x4nDB5nHlEYJIcuLL/Qk3ysigc3ul+lj6TXrRx/Ww0xUU4bupsSJXXwTBNO4EJLap4YFXLyk4
jXhbLSPYYfaZQKWuix3xTTQ6lTZ3teFQrV2CVyhJqD6OcZ12d1aaA+OAqNRmSCXKrzlhewHMO08x
dKMiml/l3q5OkHOJm4J7/NoSltaXVQb+hBtN+SlAK1lRhhvQ8hVsOZz/3zuKgepUaDhWEQgjueR6
/ypIWK7sA0FwRFJqXHfUy4JZ1MxMyJIOQ6Mmr1RrCwiG0Yaf+sa0GknCO5tSSvDp1/V0EOK8zulK
9kiyIL0Nj62vg8IqnD8LQS0LWTnPeJSnEaFMvloenPmGA4OQ7o/cIxO8ryLexOiW49JWOeK3lEco
/PDhM3CB1ebwmNboe2yVVrUwLOMOs7BDvQumpxPAwiD0q4zUAnQBtMExd2anO3312dIDyeTFjKIC
jmX65dUBLduxw/wkNRpbKivWrDkeiwmTB/lYWUdflyZCIrWfdp6tIDR0WTtud3XLH120L8YmTp9x
nQwzx83g19Hcf4XW0R9dmrFgLcA/RIYtCQlKgmIZ3yzasyhuGnBxwwL305Hfw91K6GAubCs1u7bV
JQUmCu8WGea1UcRF4xNnzC+XLIwOCSnTZojrtJ2irKEmpnKEqO6FRzmLaTmcp4tarDeHixGANKQ8
1y+0lgKx/tcohhD3snxN+15XMT+CPlpi2nv6VJmxgOst9+xEXmZhmJdDqKFibkouBwuhP227QIZP
P7xhisubtvZUUkNJwbDafrA7IgWes0p0x5IzPabSwdMQoIC8kruIx1X6TvUCXjRfCGHMMdWi3EUe
W5UybNzEUR569lj2VcpLYqYxZbznAGpQEqS/Xz7p1JVE1frvZVcDOY/N1jfuHa8ZauIlKOO5Fg/u
kkOA84NOlug0cNOSUWKF7C4qncTCyEnAeKyg+wdAWJEtempuiRfonQiU675t4Ev+53KT6HXbS6bD
qLL3zlh0HbcYKy87x9rLe1zrYhG56aOt5zolEW8lcaB/WXhSOVoSS5lG3jSTkghOGQHmNM8doLMu
knnUNKXga7eP/CCm7ju0iI/z24sIMqNoKPC42X77Eqr8e+1WGyFSTxyJbEO2H7ndznW0wQw880uS
dZQe65PQ0jjw3HFYYu8bSUOAL89g6OhURXYPs56XDNqlDiL33Z4EPViGHrFt+DdXjoaFuR8cyjSK
SRWI4Uo4Swgqj6aLFSDPw7T/+FBDW6p3Kygu8UzgXGW3IWhilLZoR3sS/DQyldukadNZXvkTcWRY
CKrRqn7DTaFnsOnAeJ4+yzSk2+y7BX5tn8A0FuWTmnQGUtfzg6+YmFFxW4rvAVg0I6kyCkRSUiSs
r99kaQEot+Oy9/4ULhTT+0YocM35Y5bVnf4rcOY/P/JR4Bc599IsjCeFtNp1sWaQH3gOXHKYoXlc
3mLLGJ4fBrw67iumL3Qv3URWjx3Xl/GK9i0NpATLHo3cwcW6g4b0ivUKC80g0yIs9qf1wybq97ab
FysGLrMEgo4b6Iu1E8nU/j3kTmlcu1+RjHamNPuKlmlKBS2VmQ7CekuKopFl2jVr4NBpZjF10Xs1
d80X3DfMQYzJoPlBGT/mMj/ywwNCZs0aTGgNPTvr1tUAGl5D4WbwDAivjtjHcQGF7hA8/G29P56Q
DKgaR2HGJd4yTGRRTSYJcGh/9oNZfxVxjoDzJ+mg0+CYEpHVAPi8EboKu2YB3otyBWOTNyX3T8YO
AEhbx7CkT8n7SNvwYsfySKDI+ybrPcZzOkzZ0EgQ4rL1NlMWFQaXClBKyT6oNZZesdPwu05qR7yY
L00xEDoBtUzMvDHeMNu8DkexN0UA9S08w3658mn1RP5ZGNY0R0mLTmO2LVvxaHxwVkw0JyMnpaxV
eYhHye183YlJ2jsS3NK9SoXBVCHugn227Dz8FlDu7aJscht/ku2Z153JpckU88brBBtpTyHwLSDp
fNH5yoB4HeCCFoS7E5wU+7IAOnFqx+t5iDfL4hwMpjmmI6bRiGgSPXi3WpWtbmPh/GmPcd3h/ovT
2IT7e+dkYaMHCu6xzL7PU3Nxc+rSt2pyOleiW16Inz5x8YV7xy6dAuwPOMe0QiRHhiQwuN2xGFrQ
J4Ck9i/fN9thvKjhZ8gw2RDuvDnVstAQ+1qsAnjAKBEKD2Z/FvgBBVghODtGMTE20nzvyHk4PcrX
CpMsZzr6KoEHZ4YyC/4yBspWZMl7eCE3jx4QuRUX3yaQ5DnMPU4oWYQVwMc3MnGhywRTFdImmb2I
bJyxfHNKTmJfQUfsNzlqpmRe6TYgtf5/huBHOSw0I3rff1N/QoGWCE+f+wnsiNOczksOzn7GyidK
XN0oWkxQCXDxgC4ACkudm9+1bANMGkXAVctK1sht2ns/Gn5Wt9+ossDHHp0gZ2uFsj96uKFqXVVV
3Rglg6jxaRnzqcksImKRhpPb/Odosav/iGDZtrs+DpvkdLEpEbrzQ4qpXH4cVhiSOnfFB5G48tZd
xIvH0VLxh5YKiktPs60uxjj+fr6yu45tfSbfPLl8r/7q6qk7xhL+QmOJyEGgP4b4Akt/f9sFJngT
hEDNcC4Dr8OvT7rnixSc7iouMUZVBWsGnePah9MC1HqEAl759gCqhhiZ/ECD7qZ1A/bJ2ged/HH6
4PmPWKt+1WU37HdqFTWLr8EeICfmGsu8lbT0vYQgJXlGjivFq4OgbQ4wlaV4tGwNjVJr7RgvSJnG
aFME1tRsPUdi1QcGKMRyzKGpzMkVTpgRiAiv2bO3/VWX8OjZCR/3p8JvizpMpU12HpXCEwYe1yjg
5OR34IWLrJfeerrQHCBR8/yI1MkPY3o/U0j9PQ97mGHJmM89WWk/geeNig0DK9xngGfr0wvSLsG8
P1MGB4tP2HoTNTY1Cif6jYMmW9/LpAyFfjIPoe1lKg7wjuRU9LBvqsWtMwAbM1cj0o5nux58kPJi
D/A+eUelHXOlW7CktCsGEPhUVYyxH3jif/XnTJPYQykJh07f+WB6c99SulXivpy2oHLFwRzJM6Cy
C5IWuAO57XSrLY1QqSV8e1Hw/4NyLSKtiwOc8CQNKnB+pyrBV7VrxIKU0AYC2foCLQ4A4y36WsF8
Mfsm5GyBtrcyHCOPO3VbgLq45SFTRW9JesTdhRKh/2mUgQbjI3D83XPG/iU53oDo3AcsrgV1Y8u7
SYY8hRhM+IeEU2UOVciDxokCf/taz/ohgui2ULGjKRkyEMo2r2BJOasPR908NB4m8ER61qc0nqIl
sPoXFcVIeiX8EvrnyPDDCnhpFdXWhbjIUaiN8C4hT9Bh0LmFW4ApUMMKYYtQZlKwTaDc0eeWDBnC
t7v6VTy8MpaZz/8MA0LWJGCXcbqCLuMt+OTlXbr0AN1ALShllQ8MJWUqlRm484qHRIYoPWWi4ws7
9ov9WZOP5XrUZPt9cMzZiswNuYbCkWrNsXJUX0RWcaqJhfQopIm7tVqCUDKEVeJdexsht/s3WBXA
BYmUpvR9PETzN44rJLdnpQVzv3D7crQc+yyrFGUFG0e4NnKQxayDs/hFH6lbylYIrp5ZAr3lgtLI
OUc6EXG4VvzMnRcRQ4ZAa677g/loVWEQF3a4eFyxGma1wiWHa7OS/UM9pV4HUrevbORZ1AcIeG+K
60AGgKQK2Gzfa0LMOZkqtElqh7jrDAskmVhCizTv9uYP7Lcgi9gTg66dOH/FoN81gMONhEGQsKrZ
siFzvpXt0fI6lEn9gufNHnDpamMo2Gk5qx21ET3hySp4/MtNgDll21g35cloThqOa0nCZf9VBQ2n
d/GT8VPhz6UHZTCSLm70w/Ee0aTsS3f5h4f5+FeWB4KVz6Iwu8tti/+ZZ9QWnL9mR9zs+rS4F3ce
tMRXfftAk1K+5jBFQNixIYBhbf6hH+b0Xo3yga3lMZ4+LobuyGIFM8bMzI++qeaGgomhqIHTBbWt
CVtnDaIoQqT9ZtFGuMoTgXQ+PbTTd9dhMJ46w0NB6CDaFTjiNTZBL/1j6kId7CCCoCwHx7d6cw5K
4D7o8S5xKBhsA5CBlZxqHH+PbCzoQreIJ9FGLkMqliUvsIR/Qoew2dKpyX7Ae1i47GlNe4jhNcq5
/78lXGAlwPUY7EfV+24vM3HSyj7uFN65HH0I6CJorvZQwZx3I3ZbQ0PG6vmf9oRBYFKjx1IlOFSe
m1QcI09tKIwWozm7Wc1b6bIDjn6vpq1iR+CZnwejn1roH/XpSiU3ECsSRW/nlF7GpPCzPEYgj7F2
uOAkmRDTBaKX4Ygz7PimDZNqhCdAv3y+gXdieCXBhl5Mlhhz7IGX7kk0/yW57X8AQI3xgaI2YMhe
LjX6dSnDhd2hQR3aFqRbKQLAabIk9i5ASedHWP+ITpn9BM4zm0H8hRemv/7uVUWPMgcu0pjgtNxa
GGMRMGaHCgalfYCYxLrCzX04VzTOmRptTdmcb57H2ANV8JbKDqDY7/yfIQpC6+niwc0AgpjX5Q1Z
d4P99cysS7eYhLSx417ZMIUGeBWEDTC68KXt7z4x59RSoXH81xs56ex0xdcFAT2zlem8uF6yhGeV
xHLvem4SHj5X6KiCRuo5R06iydHwb77nuDwH9rup4UwcwEZ1kk6iAX2P1B8ecu+JQctop334CSu5
EX+9R5EJ/9dn4e4vAm7g+pfwyp8ftu0YzEoejx995y1sWMt2hG8t+Zx6TpM1D4cnctCo//76g5Bu
JnX2tKh+nGRNw5AS5WyiAxZfeDpDVJl8sthRGQfsTfJ/douSCteGs8f/HvAasAv+atRIDdaEupIA
soYnKIHh4E68j32Dm7xjc76L9D6vu7a6E5Fv/EgYEpVrldYcJkiOAEM6JHGIavS0q1K9MQLP2yF/
9EYaTL8DH7ymSfEubAofQuJbWSRYQqYPEMkdUbkmHZcacl0vmyk5Ef1IXR09g86gvRkvj7uzDuuw
1sVKCogs+LyEFp+GLtEXDJeIySP6OjaB/WoppALQ73fHmwD8yGgDMTBDPmD2pcFglm2jK/dxX5/I
2Btb5vpQC+GgDJ0KTcb3quA8EG2DfKW2LnfTlp1Z5SA/oOnBHwsnHSyJUISFUevU74Bf4cqhcJuJ
EVNrb57Eb3UqmZNao0ZV5fH8RGw8yW5zEYmXbOXk+2JQJS9R196JmzL8ST5PmVu3E4vHkBxRltXB
5b6ebrSf2BwWt6fVkMpGQ6iYHjtmNqn06pJ50qvKy73Ru65p2KSi/nyD8fvX6TyV8G6hOvwOS4Yv
i/ODEnlzRxmyLaU/jtn0NgCUNNInW2+kb20+TGGasjd8ZNKvtPoO65TvI7DI/jkVA6tf8joi8RXG
TMuvePWEs4BbKywmIzkLNDrEe5qa9TO99o1FOKyCAds1uD2iEl3SdQ5lEBIwigZAgW0hJyOA6AyT
lbW0sLhyh8hxaZvCUQ9e51mZ8nFcUbWbNV1WBFQtOUnq0pobCE5rOClQR7QaOpOHskSr9FyjTEIb
W1apb739Wnr45KYcrc3WKqibtfNYdegx9A4Hiw6lvjY0B6r0u1dfRM2bRDLUBu8w6/aoEmVBVsQA
cbXqy7bTgFx/9dcdWUEHApR65qgKkGgp8qI2vGtdtQjh4EKcEDdPPSFz7TIQ9H2JsWWpHPXSAzV0
P5l0J+VI17bKIh0caGqKh+JpGA2ypGA7ki/3WAUc61BKYRa9rfBoat6WDwXG4B1Kb757lHTyS7la
A8gJRz/Lwfckuz9lZu2Y0P2WM+JomTOZ94QnSl1SGheedS1/fH2knCL6dJUUDTUsPZpYliiVqrDS
je1hFxRTFfPxCsA3kUpyLQX0/2LSEL9WF0C3nPSEIzow6mOivKAbmA5qDip6lX5VUv+ajx3k6R6j
gCVzdco3HojJifXHxyixaK4/+edIrT2q1xTGAbNq9YqaSx2h99iQw0fHvxsq5QOOEt5Y/ARxvr9E
FMKyFlAsuTS2L6JgdtWRQJPYMXsULCqLo0Cbmeg+GlzDiFK7qCDQFxUVeJDo0hVbjTX2BxJZS30x
7r4u3XcP9A6F6xoVFgRgTWxMiVNcYLW3hFexSN6/FK6kWrhkZoMdsmUyEmECwGZmKOig8e7b29dC
1alzhBKnxF9ya7p3yV1Bo4F8GwWnEAu+Wu2LBqChv3NO1eQXg2ko4hSzKrHOMDkldbvmBDqOa025
QrDL7v+9ljwzmgbvLKdFZcvwT45tHhC+bAHStsxM3GEXVw6VbcMyqMxCpHSdLYE3LVYQ11vrjLlG
mzrkEKtmnoNChL8N4ZRqNXqjDmuiSj/mZxxWaoOqtDxpX1Xkc6kuyOP72d+GDUWQLGFR5DtkWPSu
S/qRAl/hXbgVTiAU2G2tCaGivqD7iECqO87sCd6gskj/lpqTYigWJwE3EiO8lpfSNPcLI8dFjQQc
lrkQqjuBKTLS5nDh/EbD8dUAn6NUMxpe1PxxLHAhG7yuRs9xitPQMf8g+TvHRXRmQ3VOGAqCzrBq
lvQ0A9JhRvIMCYIqfcOneIC+glrSg7JPoh5b0VZOfrV0lScE3ZDad75qmkbDB1iLB/ThqrUtAr7N
jnAiDH8dv7y8He1fiVz5pWiv+MBVeCjJIDg2eWnfe1wbZwpqPEOgtp/bftOeuvxqrepptJ0Je5qT
Fd8gSuzG1iMC0fIaHAE6/2X+r+BfVsIxeCCu/+mAuCgkzz46SjocH84yCcu/fDCaFw7ALT7qWeOc
eLqiDAFFUG3c4CR/7bsdJVSgoh8MFuuEVJ9fEN8UkY/6RooLXw0c5lPuZ75iyZgdjsfy+S3t+5+L
kN8rtx0Uotq1kqKHOzrXLY6YEe4RNb2LP1p6mwALu/XZ9vTy5xbWGjhCz+Ayt5wi8vLAruZzx2K6
2GWBVSlIjksvqK0qwxLLdTpOBzuxPiy3XZ4ldvndUnJvNRCqmFiskHnZRV4utjhQB68vPNAtjnXQ
Cl1xoadbqds6uULeFeFfRYbZrwDec+LxIOgosUE8TWfXXZVZtbZxpOISViXB+fz0ZXXyUkTJbVOJ
qmSxCkQ9gqDGqxFOtQBZzCtZia2e6vwLKr57JFmFzEa/TDRoGPgqj6Pna0LHn+mdC4eICmjqydTS
w4G7BKfEtfyqHr99yzTLDlTH2md4OQBMwKK32S/ObRDgjc6hnwqhBqkpcM9LeIu2Z2P/AuF7xQEx
BsagTxvAp2o9TesdbISTJXSoMxmUyB6lmhU9KhyUgt/Yi0f4FaGQ6S3gR0S5OhJp8F0iXIKCrhba
3dJMCGP4N6Us2+Gu5lQjWLoW4nevfd794CXkNd6dQtbkRtcC2etrABHcsh+rKkL7UDspwaYyUY5s
eZlIMG1cn+EXjHeY9Tq4FBmkjHbThjYrkY72U0UbrJ8hZXEvffwb5NFMIx7qFpBl9ioaR1ByG3mA
a6sfedqG9caYtGbucUnJGvOwjZ7g+Y32Oc8GNo0ILZrfR+siXVJwMSRkZV1hQboWoBpJgwZnJzBS
fnf58MNAGERJUMHdJ3KZl+rna0DaYeRjXeACdDgnm45suItBw69XthzHFsT9IwYBkrdOm86rZssS
MdhuKiW1BSViQ8hwb/R7GnoWt2HijpZnalmiCAOokg3bTg9hQqgEqivXXWbZ5mokP5tmX89uxqIV
5wAwD8jpHEvL2rrBsd0YFSaqd1H7ptu7fz5ekmyI1zu4YOnT5lESwOEjVUD0CL8M424uvdCddV+g
rzb3AIX+D/Yx8t5ROeGD/oHcr/dlIZxQNkPOn4/YLdSskNG8iYxZFUECSGBc5p5AoaqXkamBLV4C
q02ATv7RonESDlWFZk2eE6E2ncrHKmNrQe4UMKXwuoosogdlk+V9n5cd4meHPLrk3/nEZ28Yyc7C
LL3DV+LJAGlVC5aOSci3FL+7Qy4sMFToPgaECfISprZBWDIL5FzjP3St/8v3FgAOlYEK03aRP/Tk
sFEpSPbTLGpC4hgFBk40jeM4xXizoDYDPegx16UFN7lAeXxv0GXH1rCxfzrvQr1QmrfJAn4FXI2J
hYSK1NLgJwXlVI2PEPUZ6fH5q7eVAOWGOQW9MEsfQvAR3NgAFpCfd7ZgJj0PgHS979ksWpCYcnbv
3Vegj1zQNKczF6j77g8/Y1omK4YXFo9wf2Ht7lNyL6Z2fRFI6CtXs0z9HFEwxzkX3VkYOApwhfTJ
zscE64gxzbPoVK36/Mre92Jir7SB6xh5ubtaV6y2Ic6OQ3+BBuxNfXbrKy0qj8lVmTFx1KqrdgQf
5iIQK0CgRr6qkhVDKOpE/EMtE+gXe/pPgL829ubmbbWXNXKJ5NfizvdFynAX9atvpld52R6XW7uS
BCIgTyrK3TLQ1Mtiq22nxs2VHf8GVA8CKdtm3OGz8u5oveTg10lUQ2gWVBR+iKmuTsMwZUUxveTr
doUtO4RIRPyj8TFdN3OHT1NrED1YMvz01iGQGxySwGDc/JcQAj4s8gUV9s1QYST89AaTK8PDILa3
R1aSZYDBh8DlkO0Bszgec3WKQuxa26hvuzqPoLDaygtlyAXSz7XG1S2Lu3VA3XdST/lRlha3hjEQ
77jsUT+G7FDWltNaUogKRS0il2lCtH9eSpFm1t0hZ0eWbHuZrrulbO3T4azd5V/uwgsfciDljLdK
ejuxLFieWrKPJKBpzfhlk980t3S+jDeKiJ6lolFrcVs5FCqXbSpvaLn+KDGMYT6KKPtF402LeRmL
SefE/yWimEyUPgWuX9GI2Sh9SKmxlvZsfWQDmpoRGKj7euPko4lJio96Eydc4cZA+PwlyWIOV5aF
vWMIKobd3gkCtSS9Aqi5NKzu7VJvK2p3KTXJLeNYBDnBE5sZjSwy0hxxauVuwhZRfTtUm2sbYQQH
7mHcoGHiQi+iQvFry4N1P0UYHe0GgI2uOSvSm3wg4Cd8c9V2WEkztJ/v+2o7C6AwwBJWAuiskmQJ
4KlrfyrB/am58iOVheJlJiu2dhq8PtMmyQGseX2Sr9ScrpS3NIkDT0TJcTFCQKwFojm+Xw91PaWs
FWXL/lWvxh1aIAn+6Xzl+h8x7Dr4QxF2ZeQcIYwfCDtHVPzOPcgnHdxO32uC4f3djma6CMQ/zM4b
cpnEK+Zn4nQQCwHNFFjUbqRm/0xteFrKXPrNH/5w1aZsraj6MUXpkmD6soA34UjLUkTtaTJA3zxp
HwRHjJO3PEB2cDnoXisuUCi4C6KVsyxm8jIqHpb9mc36zOSIBN7dgwC6anFJn8pzicfclaOAJoCo
r71qYXJWeHf4pzuhYhylVUeb6Tlo1SfZC9dWmBqiwnWK9bpk+CfZvf+4hkyqiDwyAyMYAboY2gOT
bcPOLAXTH5za7E+lUuj5y3jYNvbbzzOAnxOg66rYMAgW+J17JWF6NGEQDUxQ2VtBxJIJbYbbcJ5i
DsVS+kewHL/D0eZcYGoo1CqIFOv5TslpFAbszB0/O6WK9s+vj0BP7vymssTXMONNaJPl+Okng9is
qa3ulj60KGET3SKG0kO39zhjEXYdG2K5UYOgZrkzwcIcfk67ckTEO56Wn+njho0f+41co//YEU96
8Xo08FAyQnBg9Aqabv5ROCuv4Zf3ehCflxbwrco6Q/+4dtYyeTUE8koMiH9/Sth7caI6tSg1q2DN
9l/kpzoUMF56AjH2L+mk3oikmTOXN51ftunxFnz1+PaY4btImt9ssWBlwfJOHFx8SVwQnykkLtvZ
VIGxMRIfg7ehirNBHoJz72XROvtGmF1147ua9Jk85JQhnBySv3KRYNtiA6SnJIQuODNL93AJCdqZ
/xgcrMxzef/GE+oCKY5uDLkWsAxJ+zD1yHTL74TkXSQspmzSw1Td764ZLVZwA6RtMo+zYbZSwUsf
sMJJZF3y4g/aJjAjIlU72x2IK4+/5wOJBNvBzHoK4tQApwcHMr56A1zv8JW5ozic7oHKlhT/kLkk
gnRlDp+NDabyYcaEXWiYP3ofY+/mYzzvB2lwQc5E6eqkCB5r7sa+Jl6irUGriZ1/Ur8zji32G0jO
If62wW9VH0jx/W7Vf2Bf+Nk0bD727DCma++8nweLAUlz+Wng5R3DYql7LobMOI+tOLSmOE0EwzFK
YL0V7uvNy+GSHIfsA5lt9nhbQUecMHH95vWqvWy0B8w++9+Nja2OasdT4ZcWAo+vPUTa1fqdhdkt
J1o+nFl5V3vmN9D0nUxkhHBGJ/wdThagL2m8BqdV8OCFXpIbChWWz/UNpLcA90WtQmMoaI/6G0E8
cACtH/52o1Vo80WzyNRsEWqx6Swb56hPIfOf/U0RfBBR7jmB/OMJz9ohIOtc7oUOsRTaGMuorOb7
cuSTEd2y3ynXl8UNycp7rba23YjIEv/TRK2DEl5eZXGwp+u/mGMC6UHi+Sq6OWdbqNj+aAlGALdU
G2PBaIiea2jUghDnukMVMdl8PskcG6oNu3mlY77e7dhv8mzoUNKQu4EoZmKUmdPP71Q8PGY9FZoP
Sy5ss71CQ3DcFglRZxE3prSqlQ++Rdx8EXfPgs3BIAy6jM9VIYfnhZuCGyGF1fL3BtZEDtjMfaKt
6iaypL8fKJYm79TXwH21BI3mYo6/f7KYwQCvNg5pizyz3cVFm+jQau8Em6Xa+l1StPvuz80vjNJ4
zGhsh6LzCYD4TW0vzK3Dk+5n2dFjGNDD5swzRJbtvdbeNS5x6/YNhFd5r3kxFx1w3Rv1ENwdwWGt
zR7jlsSD44tnFoNzmwagtAO8gO6c1Pjzwemh0ngZ8QzyF+DTvUtowg+ojhyEkqNIApZUVvxE4vj5
xVPCkLdiTSu/C9TOqc4SYxscabNlmmgOE4vUqNOY8oewx2HWqI/uUq+9ZI7Yzdp21FzI0RrjCTl+
JsDEksbN+VhFaNpGZvkXbmW0muSdsk02C5OyjDJNAQBz923Lvo+xWxz21u+EO+Ri7Dd65J/3LJIk
50dAtipW0gu1b0QVmjigexACFQhhbcfqrG2bLHU7Hc8uF7oBnizHC0WHJ2an98jMucfciLizRVsl
g32QCtugI3b0Zu6IRw1SdDNq9NhXeDltJa4s0O35GwEQQebxalgDp2k4XHglA0xuHLUPrE7OxYRK
ah00ZyL07FUPOdt1yJkR1NGXJzCRIKJp2czk/fXW7/pfxOzHTMygTDmbd065IMNvscKvqRs8AkT7
oovbBIAax8BlEWABmzN6EvTIJoHlBWvZPwIJlaw+5UZ3MzuN9AqOtV9eiZ55rWmHW76AmqIe3ksr
s0yakXwQ+yHFj6ztiO7HXue5mNLkXb1/zZJZgSyLpnd03Ht67FfOAC3ZocDKZSEX/vEDVXhcQ8Rg
pseBtf8weU7pzggYgv8EOYgXGXo2l541HAZGOsOyECld7V+NRB/QcLBT6NO4JXXoxyb0d6jmvae2
Ij8Go7MVx80AWdUAvs84+Zy98zRotTZQOdUlDRzejsbDR2/UhHZyrRmNSTdcYIfJuK3mqgdIo8Ir
HYfDXNRTTs3rRRiP6ZDRmuOi+9AvOxbqKQS8iWwMmPh8Mr3LkYmWscYDtAFeBk5CLSJ0SkUJKw81
Dn5h4XVCRf6qX81srp1zvHTQFfbJ5CJXu48QKhL1JIAo0eUUdFispxj4hME4aFCxJQ8BIL144UnR
E4cNd/U5mrbWQdWrfQAGSu/j6rbFdtemoD5K+egKflM9HxQUZhEm+bCAnkO7QxctQWwYEConGwCI
MdRyZP3+7ZsNOm4i7h3UA6L2eM3Pex+5TzNg2MsYwLFzwv6BUfyYgmSkYZ068RxV5HkL0ezXI4GH
B02iCNzgN1Yj5IXkTr8Ul9sbqN7h//7kvjeZN3TciISaKtVuVDlG4xU4dXpRBdM1Mjl70YxV4KYi
7xxc/PWBFHxAZXBxvyfS2rTu7iuA7Bhrk9wmS/sQCwBmZdOY91+aTaf0S0MMNAYPpg7dkf8Shnap
MLkTsvESIizkRbErVcpgFC6ikifdOEc5EyXTZoX4kmBgfn1x6nkaRoecrO1yVrjlGz63xJRjK/pA
BIad04z7B+5onr1ELlb+A2UpEM2NNNhES3jNuHfk4eFGlb/jBvVYflEyRNQU1KsY8NOUs0VhVCuS
gAyFj6Buo2QWGG5T+uioklLqmrs/hTDnimqNJKy/rIEFJz3VpNTlvC9NWlDWUfwGw8VDJKh4edmC
NS7a8F+AwxnczdbVCiwbI0sag0LiEr3FMXHNbVOsemtE33bUhXDSk1v9BOPb86WTnk57ViqauZrs
EeLFPAqkCFKInpsFFq+GWrPyzM2qpap9ZZe0JA0vyh0Xknclmr67trHZ9cYeWFq0QTlcrDQAwgQK
ONlErdhN6CMq2jKljMtO5gQAKNqvlXsyflf1aoZKbRd9s/TprFB+AbVbWod/TA5TRAZcIZWmtm61
nkYO9U6eW0X4x0l0ABM7XU7VqPzaVWc65+JP6K+OH2ZRHZ4OFRsGTl9PIBvL4aB7XhYCQ1w7VyaL
haCWfE8eBbSBlw/PRNxP3b9om0bVmuf5QE0i/lQqERobopbqgYBgtHt52xbkjBqjU3Vesq7disdN
45ssoTsFLqq34ptlWgPFsLczLxZ/cetteOWEk+LbvOEVv/Mcr3CheSuzcT7pPqXOdw5bF9m2UIuM
9zeiCJzMaCxQTDqqsqObdpl1DxWDrMyM2gxzU7Di9ldgbGC/QDp2vC9GhkLe6+9bTtpto5GcMFkC
Wwr/Cf5KU/4EkbSVxtyBg0aExx8o8ngAn0gsDn0VM4yD6eTrTHOCtkT+/zojKywgnym6eRXj5skk
Dxijwv35o5jxfToKzeo3TQKUxL+/nw40SuI4MSzdCG+Lr5XI1wXV2lHbJAE6eD3WlztZip6nafW3
j+JpH4eRNV9KWl7bkauSIXMDy8unQvxD/NbKjvm/u4SWpzT54DQv471/N70VrdrvfBtm08lhel7Y
hDAvcq0XoBdzuAqcuBDgaAmGRRi19TLwEkxMbqk4d7FjUsFfXip/Oe9VK0B/nZi9WKZ6ddDHTikF
YwgzIZvvqxCs1blK4rZvUsmtlmErfbBuR/NQ4cZ+1CEIl6duWoOJfeoy8ZbASX5IMpsW/vLibSXE
PtGa8vk4Jr1ZacWOQL8w4NyoDcz7FhTJ2mbWmKtEMAopBuxe490meV7EKsmBPCL/ZU5brxktIwQI
o5dLs9VKBNnTsjKzkkwgiAYNMPMHv9GnWgKfJUKi3XzL3gqnqyMxWNj9OUtIfNz9tUtphdX+X1On
T1KVltTeX2uNdULs4+Pf7MOv5QAOFIUIQHS1363Ee9tyE0FBVJ9gmWIZe5ZGvs6MjygI9glBGyRm
kIlxzHzOMRJGYnlXaQI0I2JMYEyIMvKjmdOujPed7BjGpmsafbaq4GtofwPLgXm656sc7bPDnth8
cEaMh/C8fbiemaBo5fGnRVxF6/LxlTR++PW/fTx9+ZQwp8adeZWaFtANRExYWypIteWmYgK8PYdp
38O/D+S34IDhc/3/uxkHaLw2UIzI1RqD593ejT1Ba24bSnMOM4e5mZjF7aVOT3RtxW2HX+JmBVk5
Ed/LkX0ZUhRFdCbhdzZVUsgCVtqdF2rG6gDViuyo1BkxfydnI5544iiWTHFbSZn3vKglZt+MphGE
AFRBtKnjptlC/UWID01ckxqP3xepUrv0Ix3rIGU2+aS3qDdxotva4lm5becQVTl3G7pyZrfmu7gy
H+zR0EpYhS2frKysooj7iDAo7Ko+ItpEwgjJ7SBnk7DX1dJ9ub2MaSSVlfxIsqfL7JohOWkuKC6W
zPcvZITavTP+sJvPy30ntCU5iUuaS0h8ELp2Ew9JR/fe5Vf3uNjXtf1KJpQx7tvz3eq7uphRWwNF
pDZhelxNjs2Gk5x6uhQO4S9XpHrm/4Vz+EBHalLyasbo0nZsuvSIJZu8R5TFQDWDyPtF/kCXtU4K
2VZ7Qikv9EwZRNdhoV7HsEOzryAjY1ZAWGEwUEYmAJ0sG4ONBLr6JQaXaXzxX8uaBh75qLioQycG
E+bIU8AhFGK84uJ+aWPuR7Z8NKjGy+HjdpLgdzFeMHVA1oS0piK8HQ4WlhlshXfb+ThEMqOjyxOz
TWjKfqMbQQgPEe3EuXFUhb9+uNjVy9CAont1qxOB6BtTE+HF5HuzbShOEMahyInI/T/cOJ2HLo0U
/eNWWsqgNl9VumUw913PE1+Z7/KiFyVjh3pJ1PhfB412hm5qjAkzBpvJaf6Y/Rp4Q/pGuYDxmCx9
h6C55wyyc/gZsqKR7DUrfVfQAsSXw5xyVIaefy4P8EFDK8P/RcGZxWhzI2EhZZfjPjKzAK5MnSbK
CPv6xESUq8Bg5H4x4A4AGa/MNKpIIcfDO/qrPT1r3f2cVl8LMJ9SUFLt+eqdocUe+gaxlEEMDg/l
6OeT6idea0OzeJK64nFcKNA1Q/CBk020aw2j9hReKOeamT7qsgUdOuqDDXQnJ6P+33GeAOq8q64z
3oefVUDioO9uG97pyE8KN/K/xZ5GeeYrakW2gYkamam1kWmRIZ5THN84rg596TLPOp5Bw3tLkksH
0rEQb3Tlt9P4SPw9UNpFPtSmf+32eidSf4EttzRuSNEhsyT+C9P54EDIPHeOEAUMBp1a63TqJ/TP
mWQwNaCMeVISww75AjfDilidxtOl/JYUX/HYusY5wFF//OOIxDNrWJQ65xuJcFpLhvmerjvH2syl
HxGnnd7sme8P34SU8nRLUm/7Gov+Hw4pITK7+04cJFLZ3RDypSzG0ypqa7MmbjJvgvx+5c3Sj49R
I7Btb+3zeVLj4iVAwzoP/1PUOzXI6uue1OzfrMJTUQiVwAHiyF5UVAFJ+WPqy2FgczX4pimPxn6v
W1XIhozuNF4ptmFtpk8NbaQc29PGMDMa7KMUsORzDAyv+W78MdKUpE2MsXPdAYO2FSFQ9qgKkd7e
MflLLH0CgTI7H7nHOXFTwEBqTI0++/1opeNJY0vxZ1Bc+4M2ut4o62w0ey6xCk4393t+VVamM6P9
iKDRyS01fqMDeK/q2oPogIzciR2REYM/4BgpWKGxdJ174/OzoABf2Nm3JZUzN3ct1oIjAZyMBdGl
7KLUQmL3jMboY+mhD35LmpooiKIUzKjzRLlH3IXnPzXTyLlOb2vVL9UN7PUyIngWMXP3vkKNLsYa
unMYhVukskrdEswmyGjl3TIVSfdI2IxKXVwzuEtB7e/rBpMAKNDMwexoZ1Q2N/3eJMKISvf7ac2/
k1ShCpf9z3BFO4hcaFI87Depf/M/FtgDsoD6CD60+2vHMLz0ev6ER50eRjvKkbIij/X7WZNf676j
W87myXQQd9oXPoK84g4hxDWT92W8K5Cf5h8eCqfrULbXXdrwrE2rJBYBw+FrOd+fAjUC9McidJhE
f4KDWZYHZZCeiHb48m0I2M424PFZSsupJRFkDWc4AZLWjSYB2XWav+HcMl12HsUijTBuXDSQ9Ca7
STV2wtmDNVR2NgDh8w7kxmuhmIbaf5Vab6STMVWyE2iUudT715lQS30Hp80D64yU05EMN9IOPwkf
909MCL0cRnIk0xoPnxJrknTuHaAxUajaIKAOt9MVgbq8TEoGut0plXtZV4xcVtlRd1MnlvDGhqZD
hjOZbfDSyzDJBzS/xY6K06REwxuiEn/KfpA79d6yL037UdhpTAvpk/+o96z6nhVkzxsXT7bUuDoK
jG+I1pCxc7vAEGRSVNX5jx1ubWdEAcYBtTT7rGbE80gNDSg/RBP30vYvlHQddIcuiy22hlXf/XA2
/7hamF8GsV0dHm7HMZbcUAmyZf7Rek3NnHzhBRPTe76XUXudDjrVTf61ilsTSw+gPrZO2FxgBoaX
IEO8GGIMq2wIYIJGpCQc7aiptyD4j403h7DPrCWZm44XZt+VXncbYmFi9pXGjvk7XSXjImgP4JE5
LUOXX94jY13TtLHdnHvYolwQ+wj9H8dIhQVRKYYCqcSYfXb45Od+SKcbCg2ZVUox42Z0Vzh8qiJq
qge8CfSvt2nK9IrMGnx3abzWgkfcKv9+e5GS612dccpEjZu/hV5nnW8LDsP1HRCJMJ1odgEtuQ/6
5rrpzNQ3LG6BH9GCNF9mnzSIT1apOSHebL2GueRxP0ie7Kldn4Nw48VJiMv08Ll2wzWkZvTppeQx
EBp3ljaLoYyT32pwGCjdNiXjKjmjPVp0Y/x5PvK0wrg7eZQHSKqKPXXbMDVcWXbkm8WF5abz6g+N
vAmLUjLCZJCkIMn5i3q8B77LOyC4Q7BstRr9WoTdI5gXl4EnHkvjass7nqgSm+SWT4eNNTL0az0r
f4GFq8UMbwj7O/sHN7cnZaO5B/fNOxwfKrRQNd+ZrwDreO5Tpwizdf11mUHxnRF4tSAmZcpwpZI4
kzs/RQvj1twNsdB4/sqFh+0HNStA4hDEA6mKMoTN706W4JEvWp+YkJnRuXjjJJHGVbFqMSxZPFrK
5IMPsPasGz0TZFdn8D3uJNCGOkXEF2/Ur3lrI8WTi3NSGjox9hrzvZcMIAw0KJq9brQL4guDOJ6R
0M3v5l3cz4bmHxl07ip70VeEPfhEyNmBK15coi/0XZ9/7sGMtqnP6N52e3R7AnHAlgEjKyU3YYb6
iVZJ09w/XQiYQYAFYVfd/1mCCflcg1grPPAu0Cob/ylppAfcbAuJFcviXjaGhzPmN0fXsuri+Efn
S0pP7VBBscWOqX6q4moQlgXplrba22IsbozgxwNWPL+2LwJS8q2WrvBPk3Rc4KXj8rlcRkZ9SqwE
osIRSk9mkQdfUoDJ750isS5/mjabLTP2xtVrFaxEa9Sn9TNd4SQA545FavZhBnDz1bdSi9tT39xV
u8j5iiKph9jV9YiZdlKzvRf0Fb0S67SVPO3hrXx0/C65njuoIXobCrNPEEImnC//Fskr+vjTDmuY
VnhzZJ7Mz9FXt+hgWJiIrjV1DEgXD6spHajERdCQzFubIAvTEARQNPeu/0G+ZPNq/RlkVoXTvtd5
WnrisXUmUh3FGmPXzLtFAJJmFRQYpmTQwpjcKNP89jGtqR9ojqls9XHJsvf0ElwfiEY6dunOMDL5
2MJXjoQRB8Zt51GSQJ0gzXl1pkBP6mAeVCXQSTuOuccuKkW6CLgrxxAdXwFVszUZ2pDCgfA8M8TF
9heHSUSE+H4uSMBGEtk+PowTpieWTATnK1b7wx0dNxpR22RPn9SQq6vKoLjK1Z10I1qhieDvtjAf
j+dDBO3n5ZlEKYrmgmk4YwTWqa3E3zF9z0107ii4z3WnB3wHzI9y6BHLU3o2RI6+73rST6Vtdk4j
ubkAyDhdIMewkyc6tFG7WE+H93dMXB856DqkEB9eit4NsPMhWL9fD4OIg8PAVMbzKjcM45ivs1L0
5s/GsUa6ZbOxALq0GaQEi4slWk7Rez1HgOvOC64OpcFZtdYXMsxylitfY6828GgpoKKZxmgSojWL
D5HNsH3wkuuJY+S9VsUMmgHe0YqfSZiB1Ip5vgxvDKNYsLmDdI1TJY1mUw+L4NFNTyTFEfkaSeje
HQvtkZQ8ojMJI1bhUJHZTgT7L7beHYiSl5A1OfgXTQ7NTwW4hCKLMTHa9U1vSJHg4+d1Gd2PMigw
xWt9+TWv1g0wYD9kkyhKf5ZhH7paDP3dI8YlCuOUQv2LqAJhRb9T+4x8cf5b5dScXzfJhTMr623H
uNDBI6TktiEnvor3gL4oby1c/a7Pe8E9AqT4XY30rpopncRRMRpRXlKKt/YiFXkvfVADar+Tdktu
pPhrH+KFRY/cGPF6dqGG4ezArdENW0D3MhZXhPbNAZwtCsbcRWPjGwQLTcFWsb8DtuwoDApiNMnl
yhL40MYxNtlg0yT97/VpJLwwcltVhGXgRWLjU+mcdmUFs4FU2W+E1Zt7HGsJMlD05KlzKyhoiYMK
QuJjtdX8H0gPcJB9wKABiWzWKwmIWYGv/n8Vj4B83fZqcmAMZWG3itPb6oYmMx6nyNbV1pUd7hqm
pYnfQJYnbKrqcEY6nwqoyLcBRuubbHWYId4FV3Afs1KFvxsy2J5mDVP6tCe+rNRPhdD/T2jLycSK
O2MKdSAZfwv5u540ImMf191pEiOczpDX5gxsMbFvRsWGWUXyEsdo6+muUr740+2LZPLNBaQwDxKl
e8s5krxW6uA0FY85SpYMWKBITQr05m5B+hQS+qysO+RKY0ZKbvu+N/D739xxLOtNePE9P8Ef73WY
ol3Y4SyrkF85EquuvYh02GMAKpVMOUzL6na8aGWH0kfrsAeBfEudBw6DF64ee0kMdymbj/Py6Bi3
Jo1J1KAozIdYOhGpDpJgBLqybnNN0vo4M6VMgb3JtkewHzP6QKeejxcSujiowa8058M1UHxn0qjl
Kr00LE71hySQ/zDaRktqfvjQQsOY+Qt0wSYaXuCrGmAML4SsMMxX7vlO95gciybIYMcs66ZSUA0G
RAOFMSisUK9VYagzG2k/9CuYRx9+VeMUnIJvyJ91zI1pvwt4MQ9LPkKFVDrlua89SSGwWwVOv8YE
IPDIP7pzff5N0IJOqOWyBV3nNd5vZ9TNIdwniJtd+J/8tanK37b06QO1kWYJTFNC8nGyNcdzzRU7
KbljjsvS1MIjogvFG16lcLdS6ptivq8ZzUMZdVZ4RmPC8ssUIARa012C0ky1XXFQ//+hqWMk0Cgp
hqPuCWbjyX4XjD+bTMNbaOx5SkB+JWQKnWv4ZsorXJmuDIY00hpKPjdphNc4+Sc0YQFCxg/kWGTB
pU+S9CvsK6tci6n81ULg1VS8zoCD7DnbROUte5RpfMswLqPzN6r9XDv4hPQAarHyTVNU1F3AFTwG
j6i5CP2H46nnlL699QfC9ApjqWAH2lzAiB8VnS5qHV8arIkLvYlR7V2+B5tuvRjnm+7cFUtzs6Fx
Hg+SvnDQZkF3k5JPUhtrYyiWdW+T8KC5rgXI232dmm4F3PPGhjPyAdx5k2dkoabt/YSZZdwx1rTu
zgHMtaq4S7w4ltxiOGLjXMPQqONqZoiJRKbmbXCno73HDvYp7JRoTvwIQIEEyqTpBaK0+Vqnbrg8
wKCoy/hH3LvjcfgqhDDmyt8+xGEgFj5EIZjzw3P6sNBgu5idgpPZab0Oumm6T+BP+k5nK1gdVgDw
Bxu5TQ7e9kCNuImQRleXiydEVb+mSKXJcA3fVrud2tj73QqZBTo7oJx2jqVc/GB2EVUV3K5kuqM2
iaSDOnOPG0UgF1nP1MZxz/GfOibxS7nBIOCqT8d6n76FRfIthSIyPDLQw/xpP/xbK0EqZ0U5OX/g
7OKsv07HoBj1+zzz6A97XHQifrkgx/Fe0JmzVUz+V+lDkRaEMKbUXpYnze565uz2R9RJ7FDLMm2A
TH7YlLVxJW7kQYEseuHMaBRHdffcf6FlicJPlWorYFviMXpZoRb9oyDIOiyc8iQDRfPEsIv4VLp6
hMiIPzOND12ubaXOtqatsAY2cwEWvbaZeIZsk/CSD5NT1kEdTlR/ZPeohDybXhmoALoRDSUi/55V
67pcgR1m9zGS2WbC4LaJGapitByJezdrE3uoupGE0XuQMfl104nRnNL1CiKCcB6fvLKvnw9kkvZx
Z1pWwc6qtpifhhDomQM3UAbSFf1z/PeNFSJfU8JwLrqYhMztD6ExAgYPgRFgDyk0EYEIGPDTjFbb
4h2zclsHZh+2cPTtG+SOhZLQbwYszVmHOKB8f3ZZnqXsj1B0FHqd8v4UQptOyE4YOoSgx+Yhpe0U
BNr/8vco/VVVSlVDuUcc2lqKaPM/tnvXKCF3cO5y7HUZ0EIrlfvYwZsOg8uAwfJeXKfKh7AvYA+C
JM8xJVw030QaJVdjx5eetcQN47UVE0Phu99YTY0BZh7kLDWZuHL3M4BIP9qhhFKoBm8SG4Vn9yL/
RjqJmvPnAuRRpv1pu58RyVrhrMJY8fcYtrbIADNVnG1iiBQ5mmcQxapC/cqx3rBT2m5RflsrZTLh
uE4LNoplYbTNf2wEMcPirRNpQS8Gz29YIvExuroXzp4UNRj/OkWnyKjhJh4oDmNWrURQQntfZ+J/
jxXv09bceiiqreAvJZybWVj3qpf3eWFOqIyZcHbvFYG0A7IpK60159TAfySH/fkU3Szu/ZY/CkqY
skJmjhvNw2FItHMBrjZiVBCca1NMTY6eAL4j+Qm5ar7LSbpPAoDposBp7I0Xl2J2cxuwJFCTG82A
9uVOF+EfRqLx5ZbAadywiCdrDa+Ez0yFNTtpa8RmcDa2vjEYsdqwbOUxtLdDLWFMkHgVJ7UeRWLK
+l30StRpzTuGdY6z5I1iXrYkYnvosYfwr/do/J7mhMdsZNqEsdrfzF2yXEdyqUlvxePy1twJ2mmg
MNpKysj/4NF+mpkp8xNCeUg9knNb0HN1Q6LmP9PXzj0by+eBFw+F4Et/SQ58s/hpcto/SnXDkLOk
voAaMpW6DuuI5y9m0CXrlg8f8dQeP9pOUrlkGHr0jVuOasy5lQTgbZxMR6vDkigRqFcbJzp1CSjm
51aCzhlgvjkiK6VNZ3rOx6ZPeq5JQLnwhDNVF/iPJBq/C2Moj/+ANpzkTqkRuby1vxfvfGqGKL/5
538NWqPvlX+Zq3Vr/uFdhVf/xpMn/gDMRLpnJ/7eGx95ej+D5d2FsVY6Oj2YBHnacRN6C31F7b9n
V5VmB8dzyKCBHeVgF5RBJTWbB0pCJdvn12YT7O28IujHuu+nu8EW1xnpKlpBVOnoZaK2hvzxwMkk
I4pavzlG1HNU4sVFCRLjSonW2mdkNteyTb11pyAf4skqfdGV6QERT3fVTG8XUPM0voYi9BG2wp48
ph1gDBV+ZWw90gVmxrfAqUgqZCJ4IM3dvCMMVosU2pZX2ylywO7mpWAIrLx+F4bndirh8Qg/zJyu
UXcMC+tlwXtviDGniQ3HQTdrB5xADj4F0TmuRwotxwpBNRT+u1bKyfX52qA5cBHtgOkKUoPrurgL
+sySEJ3raYgEV9SZqwevPvgXsxYxYpWT2vbCZR1d3/5vx42T6zEAgGo+enqT3jVNJxX4g5YSB0F7
URQLrXQO5vOyeLRCgToxi8891GfLJeV3hUbtPICnPvmzEQgjEpILP4GkfIuIgGoEscxcq7K2LIrx
oIkf560iag4DZ2sxnlFjPwdvkl87lfCDoL6wrnabWA8vKZWxg+Myvb0UtWoW/IOmckM8wAFfcG4V
K4WNt2fxngTI8MITv0GePNy+FhDn8lKhpkC40NgFVKe4UT6MEf19eAHAcNS8jjbNkiLlVfhfooXV
dNG2+zHCWK3QNCKMpDi3Ov2Cp3XnLJ9TvsI1WGyOQ1e296oqGqd2Wo8Sr8yuq4lbq7UYheYqCO0k
7m14YVNWFeIFbyja5AAx3jeiWm8P1ybSzDKsSEiMIhuOM1/thdEBRUrCiyX9nHYyRlgPimiqsqnL
nkIlFelkmRCkC+5jo9K42WfBL0L3YbUftz5Zl7tQLpkM8isKV6bYGhmuFPswzw412DMWe6+upbDX
hgoF3Wavs1rkvWfj4B3GGwpE02LUOHz/CIMRvTnakAmTxKB2wDMlfp+3ws6KCEP8Roz4G8W5OnNl
1XCvR6113eap6Du2Eha6kSKFLiXxVQoZVndeGC/J48dBxaIbS5ffuCL2Krm8FsP9ue8eZzccrPmq
UdCF90uKD7K0isDtDlpdzFn9Pu3KcYJQjaKJGwRuHstx+/8hP1KD+x8YeihnkobGvrtqW8pQ3y5R
qrJp7f3SZHNUz6GgBXwMlr17xanBLrsEd6+QPET+L0M9BMWXjVkGIRNYD96RKxyTjp6eXT0rEAzW
pCXEqe2hAEgNSxvQeBbOeu80yX9pIRlu80yPQmOqS9spyDppl8i2Si8LsaeKaV/L/36QCk6464yg
MdkYgokucZmybwIQhEV5twLkqWquP+Ce82TCulYN57HJhbNh31N2luQUtN/D2RnB/ZlqxRBQmNeK
FuW+wNZJ5bD3CQmgZo/H8s8bLwtI/hbNk2ObipT4/vAz34yDhju5uhDBoip70fZq7n0ExkwHerve
GdwUP9bIHx7nxI1JMeMl9l2cu+J3Y5sKP2NAWpOQIIMhEALz3nS91ilyc+HtOdUc84gd1pqUV3t7
Vlif+wmSDsui3X+sh5WnBudEb6H+dw6KetnBXRnwUPH80vQFYqJq+AxllpPdTmDA6fv8bZFGHAGC
hl3lXxdJSD6SyA3MFb28Z9aWu0cyNifuP5dxszbfZnsMjO9NqtfFanAiKTXb7woYEVDchALUlEs+
QVx33ItsEa6weQGB6OsW44XoeFU2fJGf7z9pmSYvGY/4y2BHk0EzBOv4/X6VdqnUwAuoRPkzK1at
SvtUm0LB7Ktaozo3iHaiE+koufDPqjejGLVXdERu8OJzqWC5W4/5RbaOB7t8RyZD2x4L758r3TD7
Ogi16p40rLZM00hovSHSsBSq/PmtjqqUi1KoDuic+stPtkmPkWKlpUCGOCoO7jkZPqqcyBX+GOYq
qg9NlJj42gI2JdgaY5PopwEJsP8ftKmtoIj1FpBpCf0GXLTegSfjBFY4Dd1jKSOIZLXJG3/QGjxg
d/3dubeeAHbbkE3PgnCql74pYmmuoz1bTZYVxkF9AeaO3uCgFf5NO9Z2SA8PR3EVElQ+TlMvN23Y
bjL7R2w/PoThqQSe1kPcmslp2IGoOE4OkXXKxCt+24ul81aV+zDPvbCTObdQKIvC3DWxjP3Xx+ul
IxtFxLEo2aVQ4G5Cw/A0pzPtm/jGtYzcUZ39g6xn4fSE/PIm8fJyCddiGAwSKtLV+aEm4rOFpzwe
REFIMcOeffLyBTe7ZQVhWGo2v/OClhqRvepWxi1rRqEONr5rIShH6Bl85B/EX42MQajon88KERAu
qlINOBavzjtIFD3GlB0mXF9ZSMIivap0BEyf7fwsfuLOnoGafDUCwmE3jRLXN+h/Bkxm3hj1BUx/
sR7/q1yaNJDFuBjSQbm82TW9jz10BGRg+Z/umM5z5m5vCuBCZINCHgxXcCmDiPT0HKWXitemsgtL
MQo0/60q6j+vp7AWk0gbUB04xggp/1OtnK5th6soEKyypuqg8xQT2AsqNRlQxE592BnrMIQHiVta
SK2vsXVpMkAbmyfg1mPvF04Be4obolMTBvuxLgQ02CEOLk5qzxsoFiJ8Bu/UXI+benKlWBd7Zlyn
wuvvdNs6449r+9D8VUT6EmHm8hR2tqH/k7+a6PLYY9ZDv8kdlUJbLBYxZ0WPgD1M/K+Nayo7NwaB
4YRliV0LrqYYzOg5d3FpBiBCg59u7dvMFGZhvp+6a1/vyTXItjcDCYkxqdRzjipZBTVTdf0X3mlu
b8mOazU5f5g95Zl0Wa8zCCUAeLZRGZM5WtlUrDhutYazDvhC0ItrwJH41/AOjXlbvXQpEu6SQBQd
PQYhqtM/z4RPtUKLGtcHvMUPYoIFtbVFgiQIavT3RtB3a/foD+05L4U2GQj80Tq9QLqfTs78SAib
QgoyRBgYvPfAER4Ln0D6HvM9VAZZ+36CXJFtlvt2K3cj9/YmHKoAPl3RArTfoZ3iTyTCWxwldOlF
eN2ck5p6428E+piFUhPHNzEKJf8p28X3/9i4WrK7vfmjdwi+xGyVaNBFqRlNdFRyn9EkI00n9ckZ
DqHH4XIH7DGhAqvC/5eltIzJnxdxOsuM7OMGchLLJs/4UwCpMCNwKJo1rqa5Cn+Zxk259WcvjNE+
YB0RV3TikRgQDVK0sE5oI9ysIoJl7rKnVk1u8QlSxx1PCK2CNyKUDtbwW6SfL4f8absb+AOehuTS
yCszJoMJ7fsTGhaIazj3SaQWFkUMb30pvi5ArmT22WEkOEjMUWWms+HSAOXbtfIYHXp0WawOmzb2
lkBCPNfILxq2UO3M1+7LXy/BWkvssrrktL1y/RUqWMiM369tvRRTtGfYPsJLkLJzuNbkwp+lG88i
o3+bMvtzAfglnT5Xg+T/vcZYl1QRxt/wHMy4DyvD5+TrDr3dPyJcOFPh2aGBrsbWPzz7Te3bSYQP
ctUum0Xl9jPP9pICb7EyawrKHRNVmMMCT9Slo0QrJI3kzwUDX67gPRqEguhGBLBIPV7L1tlfe1fa
gaXyHaF1JKF5vYG6O+YYgrKTdclnmUpePGuMSybs6Pf0AeShwJLj4Jl/gNudVWW2e79gLrZDDSpj
/GSpRYu21QtLNf92J9i8oa45yig8u7qJb155LLmxNDRJHwqTM/krWHqLwJxfcyW0oENo36mM9nG1
NTywc92hx6adiOGZAGPLM84yqZdk6HVJY+BcpPSZ21zN8bKo4XpC1nX8k154FDdo5sRXelm+DHf3
cLg+f/we6a/0863NbLdrrf13RGIioYMEb39qlEzkPhwoCxXY2oH1HfoppL9GlZs1c84IFPp67yVl
TTZyogNo3tFwLS+Wmz2VpQd6mastdSVf4+mBMpKW9VjLakqM6WNYii/+hvmzmO7UcJuF35D6JkhF
9T7BI+tuRFI9wXVbl4RTcm5fWhOZnIU5PeQlpBVD4uPVK8KGcZofaZQCe+TWiFZ90AgqZkjQrOWJ
hdmy6s0TXGwtbatGZW5kTd1u8kTcASKaNVg0zEeWCGTJJD+TnLiEy8bCxKVEurJ4W3iitw9RYiZt
MO2R0MqEQFT8snN0w6+/0f7qWObA4uUsNiAJsWEv1yedUYu7FglQ9kDx3+xsGicKpM5nUCEx9yxx
6SM9VYe4WogdtbNZAZhEDEZZ97U5cdMfRxlAb2NFot8S2wjeJlIUKhD0L+rUqnc3dEw5EZ0ODPL5
4ME7SgzZBFcpdtRuhvP8CGe6B0rHphramXnWegAqDXcMBBEL6xjbA39KBMQVj+3klgmZuDZkd1Gr
eWm+ik9JUmR0zdLtWhqmgmqkzBbg7onVUHaMJBf0ijjJAKtsMJfvF45I1lG0Fn6Lf4Vm/PQzVP8o
wMpDSAPMLr5yTBNdBsC8r5T5q4wa7NDsC/bIBqzhMi4zkPPCEY6mHBhq5yJg1uxMu/8xV0A6rVUu
Y64i/3SK6SFpLw+SDP7xWy/9VNREc0Ifp1uStqkDD4YiIh6P71RG+8H1ss2d5SThBN405mc9+vXb
qnnvuxNLlCaMDewNBPjaw+B7QrRHdeTz71OOnDq5XbKz0wJWhRHD+mbQPijlpuVvaDUcymYhXZsS
8yKi2fru2oooapnkkuqftr/MJd5CzH2NuWFxvvCUm80Vii19eA4YmbYKRWyUvE/zvu94Lni/wQkw
BXngJxk46DA+lLM4GFf9fHSj9FkFVAtWrZRRkGZW6fN/WZPDbSi7GmfJEn9CUBa7iYq8A8C4kk2M
snv+65wr8GTBMCBLbf5GU2QldirVXvVGMLyp3apv6y3Mb4dRAn7hnsnKeDXF0hJudXn2CeJYqO1G
6VM4qc5W4Axw2H3IkeFUBiRPS7OfKmKiB3VK+gQcvXGCS8G/y6AjiSL7kqcH/nt4Nm+DDzFqK3Ao
nrZ7qUIgDKBnpyNC3l+bTmtj+y/8kkpGf1bdx2AMFgs/eQ9cjxE6QpknsrcHiikD6pnLhr3VWqEX
nI0eKhOdfwCgPDdyIrI0FR3uYT+f4Rohg2ZzumaEHNxynWdVz1R8CQxI0R/M8LSL7pRpcSwxLE4l
K/8KyIjAuPFLr/cSBti0ospEIBmeOkP2hlO59yLy2FMlTSM6EbvSsUKUNdYhzcjbS7oyh3PNHPSv
XGWzOBrUwy6urJMMmrvg4EQQyxoqLRjzOgrH4gKdkv0opsHGh/ui49BdpcJGSs8F8H1NiYG08r//
uWiyoCnr/81TxOG8iQF1heOuWVu2a1LHiC74hOXNHDyOJtX1cVKefJ6vWaX8InxpVf7AVRcwZX4l
hvPT/SuqQPpCoAEOsgAcRGTSmkNGRkXHyhSvTr222b0KYd/zS8KjcSFoAmLi73l479DStdXFeJq0
MpybrLHKZEF6UA5j+8EhMmmltxcH+YeKEHt6CpqopsgygBusRSy7Fj9Epz+G4S+a8yHkdTHP22vn
rED99pqiNl+ySnx63DBaMcNlRwvbD+c87ST/7KkvJ7au8NoHrbvy3iO4g70OXRr5rOZHoYB3km5W
+X8UiDo1o63ui5pEcTD8Y/bdmnekzKDW/g/021Cx4SNJYb+nWNbsLMjZYMcSLZb16I/Z7HsmeGLT
gNtX9Dcuoqmiax24n0df0TMAcz/H/R8COIoPBaV0cNyx7ffzBV3GCMQU3H4zp7Tbh2KbCrndOI7a
LK8KXuqlI+DxVxx4okqvWfi1vqGDQYl8JsqgjXNRitcNb8sD9fUtffSYjayuS71zjWzDm6JIdQPo
xkNG8g1HMzLRSoF5d/jwqr3EgOnx+cak+C98TEVOoQCl58k7SyzHWK26i0PASmODsndSZhqJVGte
Fj8+P83tghDxsAbZrRHm83rF0/IplEwt3owawaekWQXCEmWH9vXVKCncN6eIAyIYluR3jD71q/hK
bFr7iqX2JljfXIMleKQoPPufcpanWjVj2Bah+EPgp+ObHWZTng3Jt8PyGawLHK83CQWp2jnRvXX8
9H1SI8SelhRdmnexKNAJs6CDZzlAGbA0mqXl/fMhak44fH5h9SOWeICuOqKwXU2u+s3/cQ/5xooz
i3BwgUaZAmIkXEtz2aJCodC2ePt2yyfTPRbgW6dRrzMKD5wGkyVZPvnwYIcXJdX5HZVau6mex3G7
N6WmCyEuaeoihCC1UVcXM+Fx7+P9ZrAtfnnX+SVtZuUT59cm2yhjqJ7prqPpefc5E3zKzabFDQmT
sGFhySpfKweklpvXWUXKdluokRHRyt6xtGtYr6OHX7TN/v1WmyD1cP7ZzJF4XmIiTuBpJ5tLhelb
l2x03jEQbr89aPkpQq5LdeqXmLMcRU46cPfKyqi/Hl7XKcpUf9JpnfWa4esyI9WchIl9q3dVQOow
pttDe0ztPPay4vJItksZvRbHWcmiGcKG2Io+eAK7ner/vtxjh1WxbLNA1yok0auQzOHE6o8Rk5io
1Na267/VUId9W4yUTGRTCQba7nRFqxV/iwjEi4L6bgfSrKSBnPwZVtBInC4sYxgPNFu/T55K8nqO
7ppIq10W3R1P4tTx6YuSbKFJvy6mTKklnF0hxkix6eS0FNJ9lOlGHyM07zYViGQAhcJPs1fmAl/i
7+caD5/EM1HgnuMOSmUR+KyEFVafraYDu3LF5Zqb8rzh6lUi2G7ope+eV5Cemrg8YVePJYlZuS+J
TTxnSlHTww4jh51GoVH96PdbuUmmWSg35X/L8By9OFT37I8apJ/ERjjWaBFCAcy1BwHni/hvkiQU
ud/pxD1OFb6se4zutTo14dAxF3kwcVrTDOViUHbQMsxHQSrlI7aEP3aZHx7AHRxFEltZgfOiEAGA
kqotHYJp6qtbd1r0fqyjX6n12ae+Sg2vOllvvhI/ag07OJu13eiUx7VA64w5YEOaOhdKQLNF+icX
oJo3WzFK/Em3kIoAZCPgUUFOdTcsyYpRq2846Nvanf/d726sc8DZnERA1c73B/KXiFqqi9EIkqdL
Okdc3/HRvzjDee79aYqRFn318AbOpD6++oD7di3ZP+Dk5b8yOgGanHQvq71tap33YJ70JPB1GY5j
CbqBfGmNxiPOnNkWNJE3zdD7U+PqB6Y3yYxiTOnSYUC49s5aTs5Oatmf7fQ6j28bBmX5uJs3yxJT
aymJMp/FQRt+LPlUmnwcFDoqb6TipKw4ZcP5hLQF5p2V1qZqz57dKF5cBN+/1BcecgZ0IUAc5DmA
oY3FQ0bGwdMn1b4ASX084nk+yefcw4ROR+oWZxej3HRcRwTACvq1ncW6tFF85OACuBdQ9B5yrp0B
W3si/QuwD0ck34FKonTIJLIWbY75xpnsOi8K6MCeErlCagCJJUi27xlKgCgmQKCaDMrZzw+eBbdl
2rnB78S4Ldm/wCCXlnFkn11nhyI5nMkR1cuzCU/HYzbPUsa5U/ShvPucBQwiyCDXuBUnNbQMarCI
7BAGgv0Mk3Xm5ujYWjxnmuucBKxMxKNkeXtr1ctpwS3rpAXNeY6nSNmgm3juH0uabKoxcNnsI3hA
7KOkWQqwNPvq2zjH55AW9MZoZpZ6c8n4aDcHOqWT4CDyXxRidXVtQi4xIdhJmKF82taytEoXdgln
CSiD0Bbuzmnb7aUpt6yNJOCslkRYsEAkpKj4phHftf1kAZ1jQAYb2jNe/W1PYuMarUDhIBlKUWCV
sAjzt94mr5Jy+JCTzcbdwng6yhMfOO8le9Lktj6qFbFofMAT6TuI/sTxFdyY3begr69qZQJ2Xbiq
fKdkisppcfUzUiTibjNSveunJwXES09fc9UwJpvy7KDb7jBianBcupRRT63m/Pm18n7L+PrNAYg2
ro3HUXeZcsNANKPfwsBIYZilyknKjsYzhX8OWIZpc/UkTF68P1dSXd1YforwJoJHSbM7aX2lkbUJ
mQGWDzLpOcYT0H5p3IknLuTKUncHwHBoi3ue2XQTIzUAWfTxuFNW0vCWpYsjE4gGR1JSUnY27ctF
MpCy7rpcIF8I6btiupTWWjseuDrCQRtIu4T708fFb0vK+zTskenPX7zf5vdyEpTPP+n0zqXYblMa
3ra9TbY4ths/i/u/CCQHRo58HaTtINn+6XzGyq32tNi1cku+/zdhYFPL+19HnOq9/8aDMVEb7PXK
YLBiq72p33euh3htxPgJ9YUyeyCBrlAYQdk98J90WtBN+dIqV5yqfyJY7A8TrUVyx/3guNIfCtGd
BpZuP+l3vuLrss5ckuvupVhNrb0cZV2p/0mxLaz8XLjaZHmZQbuU8OixNnE2GjdnmfMPao+eBFXi
VPVa/j9vJ9yY+m+ye4U+aIMN8EYw3A9b4k80NholNPwCMVn1BsjynB/YYj+i/bfPKDFFKwcOX1lI
x/TCU4w/AcczB7YvSyh/oIC0qFckoyR2yYed9Mqee0zrKmQATEUplm65MGc0tE6qsEAtKU2ZgUhg
AtBiYl0SWp0n+Sn3N46I6FS4HhNacKPOH8wm49Ns5xy2yieckK7brpTOB4CGWh5H/C5kM2DQd/qj
5Sbq0jwsFyEuWqp7iVTOlkvverstn4yNlthYJuOf1PKFX6hvK3xBEomiOXF2EvEZEXzsVZy5jne5
MSVAJtojNTiy6UI/6sj/Towytf+uF9EKrlFu0KuuFEFVJr3Sr8xCWlUQoCIpE7wTHWzjFgfVD9nL
u4jyS9gChlAt8y6K2vUeWJu+zpWNFGe9LMDEb3xkjC3/xkFe3VboZPo6YU2eXmZAB+bZA/bagGJx
CkwAzSrHU+DxU+CocUNsimgxL0IZxUyOHDzdHKpXYz/J60ZL8ufeIY174LsM17GRfzKRdiwfAKX3
AoiumBRpsYfEC/5l+J7ODdcwUK7OMNqWd/8BKNAnvZTW+mlGjxAKT5OAMT2Kv58pHHFBdUGcLKN1
D7047TQ/YcKU1psblD11vr/IYtx28HHpYmO9YWN6hH5/HnqBFLsBTa3OV9AsHw76oG0w0Ok8nTcK
TAfpl17zgAMSIrG/cREK2wg/HFjKkcETno7Fj9MrN6mmf9C3gmr420Y6R3h7+DUY7JPEFNlv10Ib
6bx7SbDpXes/p0yKRymbNlgOWyKRmkcmOsaTe3t6qUg0VsFO0eVddqlgSR8hjwf8I9RpUPoH+j1H
7m9FUJQGva+PR8Vc3G2ThlbE/5rklkUS38ZFrcYgFpXP0j7n2oDFWMOqfa996nzSUNi6qw433T8M
1SZYyGkx2DpnZ3pc0xGjppKVOXK3ywfq5j7prUVmWzQyRnYstMEj98AaC1BJfAsHSw/WeekEkbxO
3pA+rJLFnwmp10rxPdBIpTeINOA/u37K/a5QNHFxgLPKsrsu+2Tz7lxkHwWHztzUdJSBm1jR+EWV
zsxb1KeZjkPIw5gKTLX64X+SpISygZqaXUP/5p5nEsOuxIHWwhyZR7zR6eilnKR++7VVLx08wdmC
tvfgm6rOj5qwY8qdXSlo5mXNPUa7jHz2q0AEFk+9el5qq144VYIz7R7K/v5Z3xOZ5B/cqo10FvoU
bhEdwueseijzn/phqmYAixQJmmx6lhuodSVsXXWJzfK090d3B62vWAIdkkYhD9EC3DbVFtu7uocT
cvqkVC+zqRMBtt4/OfN8H8oppBQzWLvJ2SypQfRpr4MWc5dn8pl10BZrzcQj8k2CF+zNIEYIkkj5
V6Z2kZbMcYqgdh3VLN4RjCmx51MjlSTU6Z7aRn4BhhJKX5a+tI1C+L3rVlyrZE0axSzuTOqYlFqu
kDN92zNt07OFDO/KiX2murC9j9tusjZU5RN2DI+GiExhF2ZFalPCAAXAvx0ppD0xU15A84hT0RbZ
1YKsvgF0r+dOvJQC2nXcIl1jHm9NSqGXurHnspoKTa8vjDzttdgz4VWk2zY0xLqsVNZVlOLVScw+
E4HCviRfIdMjdUHL9jJr0WQ8OfJER6ORKCZjYFUM118vugBEBq6hvDiPWD5m5fTn/77yFmzFa+lN
thwIjcJC0m1542yg1KzJVLBHwGD1CKjCe0l4OSYC5XG4PrDIpmxpVQwD9DDoSzxUYK/0spVQkORy
RXCkKh4GyUDMJjZh7pw1FLIf10O2veHTfGuU6dRUAkV/fooKzLWIcran16lzgAZ6WW33pBw1hk1X
lYkNcemufo6CMz6kvweglPcV+zMxci8FNITyQPIR1UjRxssJrFsjUghLi9RDd7cxXCxMh4kHZ7px
b4rbbza9suLy+yO2YDcJ4WkVPyGC5H1DJQGAqsuES4/Iy3yuOVROhvsDgaUXeyrPKqZ3/a7hcsy6
iMILTWsuzEDSMJLNOuai14uIwl25QC5Eobb0PY+mkqyQCxTy9kCJ//LStULibm+4jjCp2SYoXdqP
epW8okU/wFiXSnhUFvJyWBf2xIH60bA+QUw/KRspzH2DhwC4ylWlqSnfjquJLeEUsQUIfmzspxYf
iD8vCSEeOKjIBPYIV9/LK2sos0rdLmTrWM4VWoyqXp2rhd2u4iZHxvsTi+DYPcJ6N9PFNRZNR1oo
CeF6g0T1531/uLmDwQCAeX8vIrtCFvo0IrD+t34Ct4cFwBkCWUegjJwfaC2naBHbmGn0gfPkfH3j
/5awAOCbAXrGg5NUkRYmsVcMvgHexToPtZclvaJiRce6yhsgsRmZgQin6ToylpZpG5cs/d8j18zu
aACmLdr1HjCnVln0//cmrdY1ZvXI6zswRJWMLvqRvNCrOxBADm/ZqsNUOxy7DWRG7T1QLIROlO79
YyoV7S5JCLbS6M+LeIjGuYbH3RqJQ7rlHgCKy35wGyJ2+Llb1loWNZ6j7GLsYNkDgQ5Mq4FplviX
b9efBdlcL4I/jOMtUbkMyfaOou9RdQy38VIRZlYPJME6x92WdXcImjs5R1UmsjR29BNdUxXpFdJE
FATKakTgIAMru2D2JpIP9MdXY4XXB6io2UD8UcEawvQP8EVZOsCjTta8xAsBPqLsFu1GPm6JDNmo
nJlUiKBSyxYoze5HGa3SsQd2n1oq/S16tLGxhRAm9CmaiYhT2hz7di+CXMKVUPTPjHSSV/KU3fqy
kpAzDhws540ZYWEinymkaDeHjOsA4DpBXGerIofXo9U2vPgX0YZ/8okWcbhWnr5vL3aUJLxIERUG
P8wqDtWsaWzy3WLFml5bBpaITti0rhpKj7FUdpZjvWTkuTvyeKBi3BnKcyp+/f9fVqNLAtqAr6dX
XtkgxFpDu2vDoRu9B96OWg8SdVpvDyR+t6cW0VwvxB9VvqTdv+ccPHDpi62ihkKcqgk/g0bV6kGm
rLrKGGfSdobhY6g40N8RpwblRbOoKQ/PXhg4eObEVGcruJnmiGR/4inPLYzZ2+ekObVT9JfYFscj
5ejg7kAMsEGF6v5fBFKauL7T/mZYMxAUJ9j9WsEW3rJkTl3E3tXbx6n++/2BDJSTLE/tOBwrFEmu
ObnCTASo/fpmPJspD6V6DZtxq+8cyDf1Za+gdjrYV8fvPyXkoVCIPk/z+tFAWIqhP9yE41zurpdn
009ByuhV+4py2CbdUCNDs2rMJHnmFaUhkSXyuhXzf78CRh/vlqqg0rPphKD8WOumlROfc6MJzk3E
zl2gbl1kIQv7iXT/8Eb0JduBfHoK8/uNxJiOwd8+93+kxDgA+1gtfEjpPQrRO45SsUNkmuj5DaW2
g+jU0O5v1XIKQDl/R92pfzc+qwWXFGkwA7mNCrCLnGjbOQgof8SaET5GwnMysehg29Z8GrWeCj49
v3RXzmWNwqjWclio/wpsedrcUOsqZKNBabODZgkdMc6ocR+D/VWpjLamP/Mf6WzulIcOTJJbG9YU
UosyhxacezfAJZJr6rK2hARguyUfc41FUrGayFsxHcgaANUQ/vqUTMmQplplNw77liFLLzrnUX/G
RsCPDXUNRoNnPlJb6IEYTAK0FGji7LEPbniHDPG+QU1eHKcWfrAWWSSdiwloqmu2Stu2NPANYS9e
TrH6y7q902CSjuCuljJkxF6H/aVX4R9AYU+grALUZGppgkBqT38GkV3QEwm/FxAnYGNPmWS+dnYC
zPOu3a3fMg/IE7wogCJPfjkVChkGc3sB1pf8FxFPMSKdP6TSiB5Afb4ENeaq0hpQEv3DNoKsjyu0
8lib9uaq5V2XlT6po9oTSDh/8u4Rf9ODraUEWQS13XE8oDYlDf65fVgWJ6nOvKDaK/c1pfhsLhz5
IDcAgIEDG94HX8bO7ljw0ShZiZO3vOMhQcldxwN/VwV3f2UPy9IozARS/nhH8a85CoO/5B8L2/en
T7rvZ2cPb+RijJHmIfMHY3mKwAWtiARvgF9TTrl8/NYt2I0PVmk9vglZlHdWfAzixjh86eybIlOL
NYZRd2a8LUwxl3gwuNwO7ZjGpdPaD0RiX3nwmCdGyqzLbAFYlMzpyGIEkJcp8btX+x/6sbhBKHQY
kpqfX6OGdQJqTBrbM3JAUWkAsRuI1GUD6H57SaGM2KuO1jcZFiUQldgJmi8n3WyPbnHLWpeZImsq
bfizeA78/SafbVhElyMrKuhBn0c5iHKnirAZwwnF1k1LmDpxV6I/6pSaTWe1nzSZ+Eyhe+59ENbL
ulNNO2onmQn+mURLQHKQ/Mjs+jIsRVlY3T0saQaxskqSCSkKRe4uqbHc2NTlbuoP2iVa1bvNd4Vm
eVSyl8duL4tU9snvO5phJsD+gGhPhktQBzJwy49PyKUt/U9bAf6VC+6F8YUSuGTsNCmMV+ADJV9s
sGRQpB8unQMbpjjzWHl4uWp9sFkawbvc7hVWozELazWeFlEc7K4SDPm0R6izyyT44Tq241htcjHR
I8NOAWeB7YxkSZqVH5863SormZlV4vctzPCQr6ZwN+9I9HDqvnLRv+EtbSUgj3+juy5FwDrriXHj
EI6klUx/QT9tuepArniuXtzdZecIidjvJarlGQVhEqXoaFzvMmnGEoSzfkJG52QMYOl0xGZbCXTX
mVVNt8dWcTcuhFRYWRSk/r1azwLmmwj9oQKscplSJ+za9G28B1yftz2LCeY2ITJsoAByYSRMPDFi
96h6lxx88xQCg1kUt4kzh10AhBVXoqLovN3yr8z5IbVLuIF7musAp6La0xm5RdCmkS1FfG6ZYpIv
bnWXok2uJ6HjycXcneBZEt2IRYplUvWekdDFeAZ/74hex7YDZUA6OgbvG/L+WeuqFxtl0P3S9cZx
hKv54CNIkUQHiO+t1ZdaU6sgbkAI5WZC4+U3CQPYvTG/dHx8M5+HVcx9wnksk5es5lLhvlH2RYA1
zWObLMx2ndgj9WtS7pjtjsC5AmGJNg50tTN8NOb45QKQ5KaYu1MLeyn4MvYHWinnDmWj0ZojdblY
F+VM4sJMlabNPICyYxzdqXkH5s7nNEkXLmvdRksgn3bOgl5yIp9kqGyAhj66wtmt9my9JgKg2G0B
omlCHpUCVTO256IpdARvO8K/2lUwMr7HJtbIafhseITdYfUm+CV4vk2X/gIHsMFK0RSX17NFoN6Q
8qr8TxKZrq5OJmHFqzBlpZpug0uETupuY6N/qU9mEX0tP1xsqEArQR2F3FHBrh6P4Bn+SytxAury
+rrBhpWIeEKv9/XeqIWzbVSuogXKaPK2MVkXPJb92BjsnHZZfwWAOrbHbicP143/85QnRiSMnUH5
nG1kVcS9Ccy3SD+LR2xBOto/B57gQEjNbcqag+YfuinLhPxoEV42fKmgdilcHUid904kNMS2lYNZ
nW9nyeWaeVsBdatsjqMfXcAmIDAC9kj8SWdW4YJvY4+q/pcuHlwI811zfSvvmlcPtil6R2nEdlMA
v1bLkNrLvDHCeLcDrIhMO13ddKLzMP9zwLy3vOopaW60EVJuaizp4pMdV/KDmfsENoRnVeo31628
DyXegMu0fLtAM9/+zSTe6ZgGHFxw/kEzaNjU866Jjf7iOkx5wcxG7YesjeVMMpFPPcJ0Gv2BrNmR
YdizGxXRKrVq5gFtUXoWWuQLsJArEzdcIytw5XW/t5D/E/6nxdEfAjTm7JK2muWdXXpQXpYf0EXl
hkJdSlqpsqR358kKEE2nDd0ERvgNllPAAAOewEMBrm9tJoL67acSuf+9g9qXAoUknkpt8nm/zf7y
y+KcVGwTM68Z4e3/Q4fkKgIFTlOF+GfbkG5YldkvWD/VgKsfJK3k3RGvi/FQx6xaZyN7oQIiKP2I
QdOQxcwm0r3vCVbEGA5rqki8GPu8lytAGrss54HVDSSWMknDfVJkrXlkmfvwNBwbbXhBX6N9uSN/
VSfH8sT1X673u143Mg3JHhjf/1payFaACjar/gkw46Qy7MQS6T0EGla/3jsGlW3khIEoGceUwVWg
4eA0XQLTcihEehuAqhasZpCcUPk5cGe1GOakeSt4pEC8L5rzsZ6ASPQRF/cIDKs2G6chXXn/gOZu
S0XFLpowX1msYXevQa2ztVT4W1h8EPH3i8TIqgK6y5XcxPLquHg+7pLq67qnZcfV+I3pq9XnjYw5
QBs/B7Xv0N/g0j90wUdlP5ZmROvg10dFw7ofZzyrscsPUlimfjZZGPm4DYSpnpO6kL5tDVJ23SlM
iP2RxgD/1+jP/yEcJbKBcq4HxY4WpCvgNWRpRJpYgT1ubzaO0TkxhchHKvFrqz5Qx36KsEhczrWa
AkkzjQqzywYcXnslQyhJ2cSwScztVWnOFEoNj0jbw63K0OdCmVnPebuqQF9uCfahXHRRQQbhx9tV
sJ8BE7z7Q3j1Bhotcn+gH7b8unzYcM+CnaqMXKXRph0U4lQ1Yna1t9tUKcMDt+ah3FXpk0t86FiW
3Ybhpi2zq59xtYQuT9WpJLhvUq+aHA59vLXaf2vCAPUnc6OS06VwYskgkJB97uIymcRBB13jMyHQ
gXCClMcyK3n8C6FJ9HBhh/Xtubu8J1vU0xI5anV+jblf7+kmz5kmNrMbOUajgPOK6PabGihgkIDe
zFLtcZfxZeZMsx+WxHgs3Vd45MAlZSckU9c5LOGa8YhVsPCy7sTKaSZNj0gFcMz2ghRUscZ3Q9rs
vstL1dqmc6s1b6gJ1cf4zKxEqqjWqTIQAqzbW/fsULpsFYr6sIDP32BvML7qrpeJHD4/QcbksJwl
UKSSv/5m42fKFj7D6VrImWSkXtXrZhKlVXy9NzKsVGN77X/Usfh1G3j0DJAnVgR1PQk07504JyJH
2BgymcID8ZoADsPiQRZB7bGawBwUU676QwzUzs30YkVy2J1TQm2Jb4IeqiCSdHx7hPs6YC0713WK
5VZbIkXeWItYNYtme28h9IHa6L6go15MzFurxOjT0POrt5/NxjT0r43DyJhmnxZAFowg4A8GBxKO
ClHRJFiGlns5nEPwXDqonnhJocplqIbgnR/6y3t0i+IEIzWxssxHewhIjYEBPIG+LiUU5SBmKt1o
L+B1NxoCF1e9LcgnU8skni275LaOUgJo8N9FhY+knbgGEEGTcA7xS4UB+0l+xhVuQdSlwld+l97z
w0uKg10nvzcEprXZxyetFO21bJ9cDx6cxz70RLLnC4wwpToTYng4eQNmYN7j4RD8R2gFFCQODsdz
TGMrWqSPxcY3OAWHNCdPrNcwu6vAh9Lp//+KJdh7zXnT+2DIisADNbetWsGq508kVgY+K4Z6Ox+s
/sGBxxWv5YvLWLQ3uaEEsG2wtg2CGNK9Y4/ZzTDeoE9J5/VbR79+r+yDGzNYdrYv3NTRRWcSCcfx
Cx6pSJ+89MeSh5bGJ5MOBPTXrcz9HBZduBH+umfp+I/JUatebmRrcJg55IXpipQ7gXMX7U8ALMTW
dS+Y8VBgOoIJ8ocj9fOLiG+3lWXkzJcGEWa1wJ7VIxxyX/AQYnjPUvOyCqtVfjuSN7RJ7bZc89BI
iEsU1Y88hI3CFoCfYLoWKv49RlwQ3ZzKG9AaX55QSRvP6/HV4cW/WI1KzemJBSAd2kbYl6SaxRBJ
qI5H+/u7gV/IxmDucnogMXix4izwouI52nFjImhWFYcMdj4e/uKR3Hivy9oSMttkIYdI8CvZfH01
ywzQMktzhFUvup4CnFPaINstvVpwZ9FuQiFu8VVnO8IPEIrGY+o64kE01W+3grgaq1D2NrE72AJJ
Zq85JtRCVWFOfNrFij1eBprL3ix6yGsj3ZZKgA3RorGfaRZunW4ycNk8Lt6AscBcPpGqZ1Lyr74a
K4gD1zou6dU3kCCdNc7bYL7pXF1QKWpNG7Rhd4D4m1okACxcwZwANuFIGQ1paTJvMRJ3fmExrdgZ
cUfnaoZ9/ECo7MQCnZu3H9T5lkYCgZybw+zqlzqpDZ4mBHcouz+mF2jAyuO2ZmpooBIRA5/NHypy
KX9czN73jFE+KJfuwgneEUiLwCvh6BGawnMGyVi+kTHM/YsN7HQDnwPkYWFN5pT7ndwORf8u5LZZ
rktxsNyrHpRR+LMl4bqJFzaSm6ZNnkDVM5EABatsioKUAPV0vTIQ2AxevHffx5u4IF8242ZZmY0A
4JOa4wco9uekGvHI7aS2iqmHBYp9BX7QFSG5q+oi4xdz2oAAAelw6GeYGiDOf1SqgkOPd4dAw/+C
J1vRZCfwLL91y9oRFdy1tQ2FoVr6I942zluaP22k5tRA6g7YJTnG+bgqSWs4FUAoBPPWxzPjyuB5
baNS69BK8gYzoX+bGBH0MUgCAnuf9iGudi+Kz1KG2jxgzgedzwpK3bmIXyJ+G+e8NfQZovp3L6x4
gh1lN2JnPJ58bkshCAFfb3Ryecr/uFt5RM9y0IkCmWiNZ95H5tHFvIv062N+90lkv6cPJChbhR9l
NJZHX4JfzLOiRywyEoefz1C2kepGSwVK008t2hF9ihSq98QXEbqQns18xJ0AFfgjYx5K2lvk9T4E
/Df7MFglb4hrZJaTAn6SPgm1Rzytk4GL7xQPOXNAfp11Tmu53iNhHJTkg251UebTAJA+NJ2XwAmt
GiPzDrrfUqQ9BuqykMYzYANvmRkhzDzRA5dfMlQAS5cz9fhl9bHisKBUqyhuq4cKMxmLU5F45N2/
TCB0oE0T1q0jPou5dnmxdMEeN1RPxAJHpHnd2knyITcDbQOjy7/ovYAyTEHkQZiFR5vkrp6lJUb4
7/ozrbqXjXK5z7LCBtiwjU66c1DKdtjgQnuxB/GTwvqMKPWOvQ4E86IEQzR3ZcYyeRc4I6k/zFPu
vTcK4S65r9Th3x7DBxpQvos1MtQi5PjqaAuuePUihzGsbyCwkg+oYD6nE6NcCW5lhNhSnJr5jiOr
Q04ILo/wJ4vnwfH7lT9BpWxtidoF0wyt/wX+Kvq+GuRxPrJXi12yn/Abcb7/2R4NL0cswnWf1h70
iq2ida1SxRM+9wu92u7yTRXkNWfKmKN61alnPDLve5/c3NVaMGUFVIOedLDeFTux5o/l11X8bSmJ
EhosN5bjZRMV/PY3iAYZVddIc5bDhJH99yTutKXPmcgKA1D0lAMU1Nqqp/es635fWqfD6WLpyz77
HW9xMl90fjWh0db7unTtZy+eq53P7cG5DjQQ12evQqgy+kBq9k1a2HQcSYKZct9MzqN812HMJj84
3Y7Hx2ghx9FasSEQLyxm7XAhaW9l+39udrXHO2fruGKPyChW9QeSCNAX56x24nLYOvKvKQIUXlOk
2doJ6TaqiDQEo/xk6UBaAyC2KTRSlfPrD1nhIFgp06ZwRQL3FBJD/2H+0KeINSMEpMQubTsfb5K8
t9MbdkD48YxL3U33IDt/qGDC4Si1civb5tmj954wS8lKAOq2TYMydlIn42Kq0z/DjO8kvfL0urDL
iMHIXksQshpoCKHElbYvfe0AHV/rUkk05JRKy2MkynEpftdF9MlhuMDRZMn3wXSgOFIPb0VGeplA
+ayfNhboAV44jRNAoK9sPv4apllAG4asMrG3S6dAwupjkjxP8WIqfm1dtkLtbY/nFBWbz0U9qG1n
x2KlbM+1nVxkIgTq71YxuvuMXN4p/9uXXj7E68VwLWIQblNBtKFfwNolvjuTjW4nIOEVQUhpsUTZ
CFeg5gkVmqW8oCfG98kBr8sG2GDdiK4YS+vVWEgflsOblqkDrSTZS2ToONX34eKbhyYGwqyM3Bw7
wDP8LlchitcTOcSNJ8Rz+KYtNSNBf2NP1buDL9ZwVq7GnlylKuWwx6zQS1FoQao9n/Pu4ZiSBopz
W/g6YsLASDIRpqTfmyrEQIn4BtHQkHbZ4VbVkzly0VEbojXWoWy+GnQ5IteMXuuUvHRxrTPhzxCz
aupdTJFNXCmR8MbceXogxHYzLMLXiIHX7tMWPL/3vdyl8ZWjcBo8PTSwKfoyMXwT6UCjAoC1PDAb
HYkA1+6YMFan3HQv190KXEI0nHUp9I4XZQPP4egPxMv4DLT+iJbSIu9FAtWH/qjjm+XyeaOK2h53
O/oCls3GRwWZUxk4vzA7GxOyL6II3bn102u3bmu1i2cWIhPUzZ1j/WYkf1WeSSofGO3CPPU4lZKp
bpEDlcWYDd03Jea+u0FXbk93dpCU83QchjP63Jy3aNPa7mA+ZaLw7booTb9HqenrllqWxscLk0fX
RyLjmv3Tg8h8sMWHaK614ucUAIoubD3MLxtKL+72yWgKx6fxiRmQM3fdfd48cNRSp2UdDl2mEcJj
lfhQSHcKIQEZp2JBctNjXejqdICsF6h1XwZweShJWP0rKje7q3VoYn9zBS/Pgm4BVPXn7JGK+7G5
w9g2CzcvKJ2Jvzk6i6kPuAT+ijCzX6dFsN668k6MiYvrZFyiCq76FrsoGS/UgXCtRAIN4acJFYYR
pWNvMqSa2H5DqAQPfIZ9Ys3ZEnowAp9//3o0bbD1Z6bpWklj2+cNRamHn47lzvWQDLs3rqS/aheY
C7+j8Wx2Y880oX93Ut2/q5DxedePT/HMfyjUoCffo4SA6bx/GOoQsDnTGSb0J6kAgjpI2J+ScThx
+W2ikib/MIeQPCpt/5GXkuYjtWDkVXOfZewy1JAXkQPVx5585Xrg9f8FDtPGnuP2Z9gsMioGYB16
gG5yOUb7DpbrsmFWD2Kv9poZf1yAnhaSEt08SPhkBc9AslIUNYoYiPbM0Pl7D34Dv00aUMFJlj+Y
1YDEN1a29wja/rM/MCyo8DLgOAJST6ZB69TnmAypoIyM5Ike6+2+eU3/LmL9GbVmDg+JLCTLxjqr
6tINlyQtx1mwxL5EYyrxU+FGNi/fj+L7XC9mPF3G7VuJLIf0zsqAm884bMkTxf9cfgiqhRiyjYJy
KE9Um20UZG94Cl9WYHDH8lzPvKsaOwNiyWRJP90QAkaIKuSDo+dTwlGZFaPpG1xyxTyJ9t5sEPmn
4JeCzqeIfaVV5huVVbMrV0I7V8kvxfR4ZLgiF8CEPlBzMBs0/IATabVLaJx+bPlx89c6ut0xBkHT
Ozrr3VqbShmNPtFWWwLQI2hG7m+vwTaqGAVDdmGWK/Dxm1jzOU7x3WUX+v64mO0PszLKOM+X6wTF
peP2Jd6mxulX8lnRlV/Qc+MIp/6AJsAWxUXW2HSSLd0T31kv7fLxgtQ2lF+BtR1bWUcx6G0cOWP3
ZgkXv/8bNJy04u8f9aMaG+8ugIjoMlkHvUh2ie90w0N/hPxS5otwIvbRGHI+Nq4LKgeTcidDCD8+
OZdrH1VgoQYHNfyUfRuGcjm3BTnaSeyY0d8aawH9xI5Eg6bmgPS2bxpFq7CPVG2AWWk9FqUvG0Oz
jc/33qi29qgDULyul4+KFd+1S0lCFgN2c+x5A9E9UkfVL+Wg6NwQiHSV6fYuLQTrDkyjTK001ZDd
PtFLoZtvUqJCOTSKXav2a99+b992rTt9Gm2QHRgZFjTVfh8RpOF5DVpdp416zAvcXkFgImVIw5Em
nga3fa3WPSNXOE+hwEpEvjZ3xT8lPSueWTsB8vIyPSsCK9zmn+6E5Db12J678wE/QTVe2yGU3qEZ
vJkD/DsYSH+BESERr+6fkYhmgNTJ3YWkqRpZ45+9LdIw7pu7NFLbH4PhyGbr7mPu5IUcJsWOqxJD
t2ks9V1rfYBiKLy1Vyya0Ne84at/U0REmab+SPT6AhKK1CbMl7ixiGbO1m7HE9FUSgKSkeqptpgp
aThIBusy785nIfKxQ4PS8JnrKzLQWLq0ufeeoVlEfbQG9avCGILaarQ5FDL6zFWAZ9yPYvFk7WLB
sSPaqNw3WXl8JycHvQyls7cvg4IWV/tNtBv9E8A3ts8Bgh0NyFYdb+yOI5IPA7TFD+0d2N1dYs8Y
FRG0OGO2cVayQDu0rWdOk8DX8IKknJUpejAZphv8q8+1Rl8e3QcpdUjSOnjVJlGa9XVSY9RfCFDk
IoiK54bmXIMsUebe+R7GfHeujbaE0dwJsIlDA6rp8Rl0hUnjuflu0qRRpo0CzkZiAGIL4N6QDMIQ
4KcxcMBOVbGkeagLg42KKIqhSkapSeG3vum8eO99P7oGO6bMGnt/k+7qsbPS6+g1JO5x691/pOnn
E8zOj0exG8LST3kdWPXYlDPoMYfsU/m2zvuknZqDSd+BzeKA3oJRyRdMBvBmjTPoNy3+H7dmBb2b
OVIxTNQ4exjX3IQJIqJv27Kq4RxUDK+QZsnPoNFpOhf1vAP2T7bH1w08VXQfvHBfuEPHjeK7XYFg
cSVi7oLzt40iP+sMz7OT3I+O6u6WMas6Sc1FTsAEElM6nKhV7nIba4WoKEersGlDW/sIOBjsGV4Z
T8ajIxc6+l9TX/fNbJcEpYlEYkzmW+X/vzNI5lLvW0pbQs4SKgpmeRVoPBtj7J/o3FuDdWebjhTJ
h0IV2DiiNWb6MUjOnzBJgFQv3DS4imTQFVO//1akjiJVsa+dn861uIjPGP4wSL2tusfphfqTkIrW
54coyVnQS1uJtzG0i9ZT7XEBPX+3S3eziEse3kNjPdyf8KC+XTMFtgM/sKFsZf3tXbDGYBs7Xg+M
iVznJKuE9Cnii993CbFVcCM/wsAneHxqz4yxp4PJdeXpTiJpKXWRarcKANPBdKMfrq+dYJNZZvxN
B2BMxckwCqEZsvd6EMWdZWmmiectYq7Vo3sAimrMRieBTgPf4EFAQOWWALQOTwVZ/FVL97e25yK7
IUZdFl1QK7KFFy8rCuklL1dAu/6ZNmDjTXN757cpYwuBhxLgQ1oHOMcnD4gCWbH0RQucIQpJRB2s
qnP+0U4+lgfijX0/0LxOlhVljVJltxRsC3hXpC5u6+upyANF+XaVKvlmodrOrL5enS/MitOn4Aq4
BaVC2j8FmiKL3Cm3gipDXfd8kmfxXtGH7okZGpgh5gi1R0TsEAsEt/+nUmI8doGJB7K1JKQJ2sus
Xyh6X6UDoC9abR0AahOuefdhy8FotL+DzqBL3beUg3TlmLVl1DmtXFZMmBCTGAGeY4F3Zx7d3zUv
kDsmShbsb+HW16fAXPEMPZ6uNRG3TYTVYWI7nB9n6kES5T40ReNm3zLWi0kbKX5VpJw5CMPna6Ms
zrq7kg/ZUXZIGuF/jFHPn/HOs3DCq1QFDbcKdS7KN4MF3rU7sBI7hN8R7kAzqxJ5CFB83WZyHNdC
44TPUP08JPXXmbwIq2K+0JCYMlTOrRHgBnnM4e5lnl89cmobK3cepAZbukmqYgJL94a5HpegbYWR
gbfZgALL4GwIqmW5uztHrjhIrjb92UWuTcSYHwSdV72CM2c0TrMZvd8GxzLRjYB8pBVRbZlUS64V
8Ae9dC+bH4q64wGgFBj/QkuJvNmd5muJo8rbvs532Mn1+ZYpEe9T0mdQZpZvx6iN80DyLRAOQpEv
eYnPTDRlk3SiSWfuucaSFC0wHJvjHPiNDIC30byI9xkTlD2Th6G3Vh8Gvoy5mUKtQaB0/DAPWaAk
7E7o6xhL2OpRINqXbzh5c8CdFbb8wAiC1S+mF0k1BCKTRkhbD5odX+a/QZTHvmrSjTlo/wcEwHov
Vw19MJO7OT6jJSXv71FKziaoIN7k0jhruIi8z4BrL7lxFAgVut9I40yedywvskgHb7fFIryvX5U0
DlUkOUvFVMuTbYSfYMCorZxCFR10spEv3DHgKrdNVSUOrtjFo7BL1lWlLUCiIQNtijI2fZrMWGf5
FA0nd/kM1+PMWr/B3agyuTRtkJetdolmKeanCmGWirs/6scjTJr6Di7/cIaeGHnNCnjS5sm5Zs3k
NhxQsBZMTiKEc/db7hUDq3WC0WC0gShtdMXGjkWgTOngegPS3Fjxu5OIrdW8sU2xbkux75wT/Avv
vdzUTCGT9WQ1oydKVQZUYv4ahJ+mamojJdRune9crQIR037QqyAOSb/FhBiqP2ro0DPRAdW9hXL2
mH3iAI6ZPXlHTX7lSUnqu9gPZGCOnh+S+UE1ERsq2IhiBDILSEdj/oOwCMug068nUfwH+1bjAZsP
eXJJF8IcilN+WDDVzKa5YOM0bXRhNfLDtatY5InVc+15D5H+LG+D84RtAvq2gXVJYmBdExsrAdSW
oYNSxYWgQFMqrB72upP2RUs/a0QSeJSiPSARZHcCk9Ji/YYz38cnE/GSULaLQfp0Gu6cLfFs0Uc0
Z2WLHktNFy98IJD+/zUPjYKMYYpjaZT+e08FoO0lZ7TpIc4IlSJ41oNmRyP5i0AsMaX+cQsLEiVo
BXm4Zkb0iqfRMwnJ+OAup21qA1ziamMjAJUEo7idZ3WKfEeCKpBlti2eE5ur5RMDHufmvIBG9GAk
bCta8KYTPo/mtyCv9bu3OoBc2+5PUIur1MqRHkqMq820NIUb+PLlnadhFpTThkmeZL0sZIwRwiW0
2cBnlieQaCYz/+By2Wzpn/ncSqgha53t1faRg88ZMgc1VuPoCd4ECnw41Q5I+eupgZimZ/iCUszd
fPEth7NyIWFogpyqOMAr3umhhTt0k2f9PYiq18PI7rUyQDECLfJJRLFIkkLzVMLqjZ3Om0EQLfCE
YIfb/Umc8kVi/18qy5q0NBwNnEdGoEPKXCg0vSgXOMtXEDWFtK0pOBIa+cgSiZGkYwfNTmKVeLYw
DsGU0GB7Bkj2rmHjM45Ok6ryBEI6yLc4LMwujsAncTrtngn7r5lOkALo7JKp72QTloFTWCMS3D+W
U3SWFHY9bI5XzZD+RRcBUEQiKNjtgIVROB+FJXIVFN2Z8HPHc2NR02VNHjWmwysMupo0No0U8gYw
YodMjR2A6F1oxpw+UwFQYZDxqZakoWq9sX7dLzrRTaNKUkNWHs2yhQH1y9lLLv/Z5W1r4xtUjZcj
4mc7l3+/wTovfWb0EMCKuIvxr5iRdC105bNicsc9kgUOFtoJ8LZNtdgd/acSoka0Ov1AN87lOt6P
CB7wHOkeC5E8TnTCwLsVqLusV+ANl1RsDKnXiOIhbLv8FCcWvUVNtY8RMGOMt74AFPhLWssqfBZ6
0gPT8o4iM/qvQFQCeWQHdZMqwKm0rBtbC+G+m1fZ4OYPG1SZnfcBV9JrQbhhmBY8l0p4LxOcdqTV
DwNepZiDbYTB/dawFEdGQtEcJX5PLzelJLvLVt7F7uagU+y1O7N+xS3XvG+R+wsdnLP97W7p6hkS
g4SesRgFYaUHpsJBe4P+h2+0ejeG6XeUgDl/1zBINM+GoIEw995a4vRldjkzr+Omtr02BPlwO8Iz
fBJkSgm1NzqLaH0/7tiiTKABIQYAZXxXDVpot0/+Kp9kBF8sF/PwYr2FbYSph7M/s5bsRLJoYxm9
t/iC9OgTdyo49uUSCqERf5n80xEBI7kzKTSdX/3u2y+XYSllH/+mOwQf5Tjdg4Nw9yzfS8+2aoSb
P8jT3LB4gqQIqt4poqhryyCMJgeCdjL1C81RptjK036pd9mYqItKNHRFZ5GmrolCZkJdWmPyRkSh
wdIzJ9mTWhFT0ySZ/V6ZgJXmrkAK6WBNLdcYKPKpWyr6NXzGLkiOyuXJUY8XZziN9zWMiYyvUu8U
UL3UhX/7CV8KjqEg4zeIWTXMlzZa59clFrzgJwLc8KvEDtNZgofcsU9A0aqC/50jR1I/3Tel1GaK
B/CEq+S2lG9SJqUw6d3qkeyT95aYAfoqY8W4q9qzbvqSVaOuenK4sUBWaPElum2AIbh+r0KCRmvN
yf2UsO2dYropsw0mFI8pXOPPNM63FmEzA46cyd3Buvxyb7vQ13sffEBn/IM5qXyNJvVT60OlE0vB
MkKDhrHuZ1406zARqde6qf9WFPHRTzR3wdeI/qDOxZZ3CKIjJK7iimx+pBQUXPPEQ1OXEtsopJcZ
VmRoXpkv5O5KBEODutNr+SxjsdyJuY0T4PV1CHMqe1XrcygXhp6kA1QexcWhi6T/cUzOOz9LuNuv
mjEtnX3qK7krgu0cGI30R7v1DQfF2O3NpuXjJ1zXq+oBvxfkLOWYtGjJ4bDM3aoUtPmOneHpGlbf
NPv36qAXleoXCtm43fOrpI5RT1MNlnKzNmu+ZFgCH7eqf+ScSthkSoSWR4DnQAvjQg0JBy2xashp
G4MtOwHOLZvMgle52kWZg6LcBBAmhcJstS1wbxf7v+eWjYRO+KGnphbCtQyG2uDS45bdqbHK6QkC
EflsayUr66t2Jb1SUKunbQ3IERSnXWoOzeJKkliNI85YL6Ps9yJaO35BALoAH/jGB+oW1DS1/XH5
dUM8zR217UXM9mRuR4AHtW/GEFvQKSP0l+2JkYUdMSnXbANT4zA6r2I9zBXqRuChJ/fde5f7A8+7
cMH3oDDy1VeHyrqxd2WEdmDfNn7tap3/4WysA4Y9A2oeeEoyGwVmItpAws7cnW4Zu8VHlDJapuDC
bw7gi3p7+qCHCNhH+hGghabK5RkCgHaE4qpsqzW98C/mOYkSpCbm1dbnuyNVXyzBSE9hnILgccU0
OILqMoGS2AHf2Yqa3deTYq4mWOun4NBELUhHJwNHITivaaEbTMWniNngLS3bPJzcORlKsXLPVh8p
HLfPadNXJJgY+udxu6A3kDpt5nCLp+NOwqhMLpp5zHuJ4nWM+vZWS1wzSMxrbZnFCyB3MZxhODok
JreZpCjFQeAyMflgoibaDyl2z97Ohir6VAUoz9XUiAbNKkVMuFRJPvlQiXTETR/ojZ98ByFtpeOA
JpzlJmVFBvVAGmZkTYPPOaKb5SpLw+yCLdxpDadsNjI9OEVXwn7cf+55ooF///hQunsKK5/dfevE
NXJbv4iqF4Pbd6LaqhcJRr6hoATcUpu3h4sndDSxVIo5ztBDBO4vSfDaA/PihK/bCpaKbBaOl8XG
IwBDbh2zOBR9PBltY1z/d2fp7eI3tjJdajs0hD4mf3HAbd0wLeIjI4BoDV0zZtPpl4EPG1l+/Az+
55fvwdMvdfmRdZghanlj6LEUfHJr810910Jmr2FvpWXsTIdJjMMN9XSU+Gwl3wcsCPmHM6mw6NMA
6HLAltBgK1zwbmK1o1ieQEqfMPmYiRHUaiL5QDZaqS8GmaH5b5UR+OoAbNbpAdJZgNjS/M/GfT0V
xYnIdhzZKm6Q9PMxscTMIPVXFLM6xy8ixMwHrgT1MhqF3D2ikHLbsDnwxxMeaVV5ALRPhsuJPKTl
kVoeP5P824j7dzxDtRmDg5Hldn9s1fkvF2HbipiC/6RS+i/B14orEfMfRkD/bSU/OLSdbumOS+BH
su/D/mFv5f9id8yOC2fNb8hC4iDinaf0QD3jZxBBQUxLjb3tRwfGZApHsSFZuGsAsiofAkaLQP+A
bd19HQ4a+U+QpSAWthT6NfJxdDIVafmx4k+lgfjxkvEyCBJb53vn0qvCSRkq89Lw/o0EU3X8MwvR
IPEWJghfDfr00fcgh140MOjNjLDK6uYcMQp5yYBXHDwU9b4C8EjX7yX4yraVhYwkals1/g5neOyb
eCeLFm4PIO1DfZGK0BADHnZNcS/f/ViYbYreH/RCH7ryo49kBTmDqx/s1VB4/9zSI3ZxxHU1bdWu
EPIVmVdFI6QQ9sz463dCwy0051DAC6X0XkYhioTE/YARzVFouYn8CLia5tT5YpOzgIRbtq6K8baZ
nT1iGkonQRu+05+UyQPpZC5uKnzz24oMHvvUNFTl/B1czdOP678UCMPLRhWpADfwlUFJd//4J6U2
wjeoA2QM4a+GMWKTBMXcckqPWydyNtFoFl/ozOl2wrC4FuuQs7YCXws+RTKzb8oYN7qwfaCJhD2I
db/8YfE8aWwU4B8Pzt1E5BU/JDsSpdg2reQrg4jQhO8dxuWoBQ66eQwm7yVrFTGv58TmYVOn4o0I
D1VjOdFUxE+4l1ICybPBMt9g1oXoLxNNGmUHctRYBiXDTICmJt5TQzoYOEwWg2LZcSlzWL3vnZZ9
7RFbz8K7iOFgNYaatImva84F5xIdRkByQBkJWLfZknczKHkVHX+uE3vo1rgPgt4RNFQonvzUSAJ0
6oTjzz9EAgD74KbnClpiXerxccY/JJkzjSWc1eQrQQN6IzBSiBCTvfZW53u5bk9sDu/YczXDu+M6
zCHn6q20lfFRzi6wF7P4ZfkW5k0cRaQa/wrL2FULsLzWLeHA7fSlB07qVoEQWo1eEYU28FbtbK0a
eA72U9yH0P8lqxrbX7DV0rS54bXhBBa416uuZEUFZJHSHamCEs++iNjq3z6vSgClTNv3N2DOIMDP
wv7gqKyA0vHEn8/5+uxzmTWw/7BF0DSPTWxXOGTxb47qDqXqTH+4EEDHjIsedN+uDxlczLE7CSGd
cix4Z8vzEd3f58KtDesVO7P4giNcSLI4LK84GEFqydu6qxrqYMklf1KWAAOMaFpHKYlyk4wu7LRF
oeOhN0+GwbmsLvyTXlOH3u3gvAcM2hU2RG1JWgQ3cJs+/p2FVs+jsswBanlGvPHaoV+XFbPlnF8t
tcgQ33h/7sEyHFp/xVZzJwvTYXmcPN8Fq5bFmbT4Fas6MK4ql9G2L0YNme9YXzUs11QHLNvw63af
HOO4UeM8h5X5zYcrrjVPSyr9MOltrjpvIJ3Js/Ce/VjAOd+kRI/gug4OqixcC2tm8+4EPO9jWJii
47Eqcgms32Ajje1oRD3+8DS3lFRLmYHa21qu1YqyGv4mjd0k4yUzctGv4xTXqFx8ILg5c6vdq1K3
UUgLycWh27t6cUabtwI0B6RN1t2LiJLcUxNXNP3SBL/sRs2nf6SWhPK43kOGONIvE7RLAGMlNEl/
knA37WCIKme2WOKr1BKqazvXLOSxqeidZnsqLuMZGmOOkP6AC9p22IwxuPt146WFRC1l8vb4qiDd
Q+KQ8cv6mUe7DPb3j8ImbfnRZSwuG0DRZRvw2m1AggpldHiqF49cZb2GlAkpF0urzna7W1uSixAB
frL1d2miQJUE916qMBi7uLOjbdzkVMrgRr+9RNWT+9k9lH6zIfYoiysLo7Fpm+nX8m8rJ4DkoRpA
ul0VyYA+doAO0il88WCUYjYJYrUscwGS5MNYnlmzamwzp/uZf0Eg4p2YdagPRpPl8A7Ugk+wQQ42
u7n1br1hFqH4Y+pismi4N3AI3EQu1I9/UBTm7IB10t2NdmGI+yqFoXGP3B7Zf56YWp7EhbLtZXUQ
ARYFE2l75oF3LGD94o/bXNgZ048d+r4hOWYydxUiM/9bMmKHhqVzdB3tpB/F19+ca3S3gJbog0GN
cTMwsiezvVlEl0A5PNQsMgziZoot3/OciyaEJDXQ/046F/tJwwCULDp4mQPtf2EDS1JzZi/Mt6ha
yIMgrbJiUshyAw3d1z2/s3SAs/2NOU1s093huSgottBWYqRFn+QgVXaCAZ2BbKIUAmvqSCyKS+vU
VdZWWpja3S28kP8sgtBkIzn46jke1FDRz1AIjcZ/VnPpFR/Z5bkZ5COWtvxm3lzhEL8snpje6vJB
9GqJrb+FFmHZIQjhZn5tX1m14LXlhhqchIZYQGTIly+xKFH0Pbu/NILPA5bE2/SLwbhYwK5Qefzs
TOU2AFB+6vjtZ99kfUFIzblajRwo6iNT/6c3cVgMDQ7V9T6qOzStmk28IAf3Pyvib4U7xZ3CkNui
VjwJlMCZQkrVSBip9pvVtBoohSL+tKncYvFkmQmtkMU09J8DpdXdFJO8D1M8gNfRoNqIf7aYsALr
cvwXXzNj7kAn6Xn9oe4ZYRqWkk9A9bfSuPgyXMWADrqTOVqEv1N0vpMCXk/RXzTOJ0NQCKkeviNM
iE78yoHz0iCz4rD/0MkebiyAViD8JQtS+02/7e8h+OODyr1dcbd77pXEuwTIdlc4a99fgcfwHssr
JQfiAhj6A41gU3TP8af16a1YP9GmWPbuGzMo0rZcIAGHmZfBT4u6Y9T/J4GklZI/h1k2KzGk+LG2
h/wlz2WlmnKvtP5hEM7c1AC0PuxX2gJm5WiDOSWnG8h/JVUc7TRYmQ6rfXlqdlTdd6AdOKGkQEIn
Bvwg6dp93tLoevug+5y/aCOQqcNEhZIGYRDSQjcrP/i8ZyPzbqVPgFS7osjXgeaYxDa/0/FzgM9P
y/LQMUTkk3BF1r86s8qio4N/B83pBYKTCXbu7u4em4Zb2gyx1cQYbEEw2rOduWDJexOx0CG2sOuF
ZWl/Luv4W8KHczY5oTWvTuLbQ8gFyMKDQ7kM5PArnwDclnu8yUUEAzTBqy1GN+iDEhsyHEbhoNY4
xbhfR+9HoQsZB0KgLw7he6nOTAPVgNYA4l3iRTIWuF0QYnaHy+8pHiNTmDLQzRsEMFlc9MsQZjIb
j+h/1A2ugT+yFQjvb+bxHe6r+rttXTYlmxgKd0d0lrQ1eqN1EfaWDPJSjRMBm3OrXSUHA9u5sf1L
A5Akuivf9ayLO/0j0wMqevrA5YzE57D0CxuyavZ9AUpBJTvjhqa/scaNtrte7C9MnmhFQoO2eyV+
6GcHGzNbUJDXmf7oczjK7oJ3rTeCq80t1CmkOXizpGy9tPUecJbaaFhC2PO1Q/64OvcZx3FTe3EG
n1sO0kQRF42XreNw1eHnNuE4Y3sebN8UiIcKMbAuN5h1mhYTrExUK36czOVNSaf1ZaLDOe0F0UE8
VpfCNvSP0Bi0LOgBTPbKpfZllAR/fD0M56NZoLCJluRY9fU+R/MjC4aP0Kl/l7FhDkYCuU2UQgsV
/mlTIYqMeDrBd8rlsEZWxSsWyolOzQ+WgChcih6Eg3SJ4AhKI2WORe2SmDdxMHRiYgpOxmeSjTo2
NzwAM6XieAdRBRdT0I+Sn/DsK7tEqJSBlAXHGWPkBszG8MSgUFZNHkZRGi4rwsPjo4i5JClQV4x8
uUsiLTmgwW034Xm28CE3BDW3KS6QtTR8aLy51mf2zABTe7NkDSs2w38UG+Y/J12l6AvPHGUHBTBc
twTuTUou5y0Hm75RT7xmQtt5jYc08LgEZQOxmryPxSQ5JxG/4EEaF35EZlSoGhhJTM/K/+u3A/Pw
LszrIirEK40X/rcCfcX9ZggqHYoB3XaLqPH2GtgQtNBBkMc6xeSHaRPggGMxP3eP5xyqTXAiyQq7
B/Ocxbr2C3/3s4bSXB8LuNn2T0yyjO2QYkQGwYu/sk+8MaWMw6cw3Z8BCSOjyXZejle6Rgbp0Cde
6Q3OMsyjR1yZUXuwFPEv0dR/OWcAsazVPi9QVyqLMqrHMfjv1xVYvN+Bu0C9ez2JdHCUrfgUL57e
LvuHec7KOpdzrZ9QrRDIUZMQLeCad449qH+Z3ckJo8NgLEoioMrlzKflhWuzzkTnSHwB93pRnWIi
sHeo3j8qG/wk8nAZEZiZJe2NYsVdmoLdtcZQBRYMkJNbf7GsXBRUSod2GnB8a9du97iS1m5UUAwq
B4FIy+9GDPwg0YBQRnye82ba5M5eBbcKA8CCUyjcf/ukdflN0n9S+Z4ybVwKFIoFY3BbOOle1ZB0
M8Hgni35TRXgh2228L6r8p/2kq6SsxXJjlfsAVDlbjTXmDvPiebGeKpaLAJLfqPUYzNQ5O2CVDaO
W4HG55zBCxOmSYonqv6OXfj7t13upnzKSafeRkEFvVtYZJmQLMfgZVQ17yQYMtan9gadA+KIwCEO
7u6dRYz8rKNsnE+bhtJs7Iv659Zezuz7GLCsDcVHqAmjpYIx/u4We/i2qsAglpy8ZVSfJO7TP25V
JrmzSnUu5nUSqSSzF3Ua7SVc9vkaZdGM8kZ9JmFkCwH9jRnCu5pmQWjkWMh083aqdKKUR66Ce3rk
fgy5EsgLuQVexWWktnYVOhYziQ+NikgYBQzIDECfClXfL8u05i/Td15zWyp4V7XIMkjYJoVBn1aq
8gwpKDEiHiE/gxVCPq8AsLc7t01fxigABJKLGQAwRyVPK5jk12JubD0O/c4WScBpvCa0Zx1Ekoc8
mtB5ggeSBgWx/VsXSmlZizAW+rsgro8Eg97ewVJl2lR+NvD3HhUpntc/cLAsNf/N/NnUB/6IxWZa
MWLzc/+u7SKqzVTFJURWLu+g2Tdu8GBsyfYA5l6br2O0QmY7pa80mXJPGPBlLDMvrtL+MvmrUW3F
C8wiyJ9twIk/+tXA8fBQ+YB1LcavxX7a4nKIyfYFZVkT15WPv6IJPPaHrve5P5DlZShR4K3Tg+k5
W6MDRoYgDhX6q6TpaRyRscWKV6KJJzeB2LmGIX+Xn89aC6gQVy0hDvoIxigiRk2+jFWL38cAOhpa
A4zmDQJi1Pe1XluWLy5WuQtprxVsspiG7786LwdJu9Fle16Z4EDjIgaANMubz1Cusqy+3XFwxFeb
tXKYPG6LmOar6jFDtMDPA94ILJW/oX+xkMfeomk8YJyNrtsqOi/lo2e3Atc43lrvcMhWubUuD/0f
i20MjmUVWa42AkBHZdnDjx1nAWMC98nJ/1ic+MJVxh4Ad6SvsmZos4nLZc6u8xCLJbnQPbh14kYL
4aV5nChhSnxgR5dQtU65k3KjM+HWrO9wtvpl13klGNfOXcZsn1srdPu5gE+MY/8J5ch1iBg35R1x
gBGIwbx+eQYURaYGW+xgiN7pZjDQesj5bHMdFvFsGYQdINEs8HQNrvxAlNrchwW2bY3a/jcl6ALg
V0/xqlfVXDapNOqexfreTji8q9hN1eHIIlEhswkbmMQuHJL8WMHxC+wy/+5G66mXQY8IOdkfJAPr
NLAiDRSGcZq/1EniTDoNN+EMR89oFoxS5h6kCPdMJwMr3kW7b2/3RbmdPLAVpPKNRpikonTrm6Rd
NAK/idhlPEDSvYOSRhPVJHorSx3bd+MMrK0mFMv+Axjs90GzmDOQipYqrI6jUn/ENgC8jY0bksFy
GxFDgXlRjaca/h0BGJzFNF/+ao05vTByoME9OdBW+Mo+wyg8vNQCgj71UQPtbisnWNki8LjcCO1m
Mn2k06VqXSxQUzMhbwWurTZcPGgE9kE4y1qtDpiE01hSANYOGlw0yQ30ufsGeuTQwCPsmgk6p8el
tZUO1HUNVagNmTx5NWIOCwth0oNbAMuwiql7vUCMKb6QTVWPcUwgFLS1ac6SDonpmgXy+7xDqgJN
P4LJCBh51oSSvpf85K4f6p8lgBj36/h0laMZe10mdAtEpEiyWuWzZvUOkt2HR7lYK5yhay1G46zl
GHyBR2xWrXj0QnF+4a1Y2xkcz9GNPGJgkTTNAc5yvl1fANckSQ5HS40TjkQeHOECOgH3nnwGOB8s
2nZb/z/XMhuHq6+dqnpKp2+4k/EPlaa3HMUp/vP/k23XKIbSk0G6LWNjx60DYBWCE3t79qIK/TnI
7K6HPcYhdhUMtF2LH7+Y0Et0KPgcgrQ8BSd+ErOzY3lNiSKBWACsj836EPJGJFoMauDoITYbeGss
m9VEwHP5jqDsKSGYOo3yuXpw76ustpWiaQrUNj7rqcNM59wALkAUkvoQijPyRgY8oeGZA12ABLrv
UaM5zeMomC0yu+qhkNUFzB5TdUWUMQ6f4Lf5C6h1c3rMwHAuT3tnBOgU6cKYs8SSGRJf9mvqMpNf
lUNc3eDiNWCa69LItV23mZhw7hZJm3poPmEzFpIddJltqg55mkzjqaphrbNMTe21MJpncRptWW1g
Aeqa9uXrDFo6JFQj+z/pFez68azgpAkYbQjoaCLL+qHuAhZL1KAvQdg4fQnLyS68fEs59pXl44+s
XhRs0HrS5IR1Kv2GOZYOFHd10JHWBhvvmV55qEPABqSJV8CPazghb1NqM0F9XlUmOQDCrhyuh6fI
lX/TSgzNAHU0vPuiNSaIwLE9S1bDi+naaqEjSD0sg4Xq4BVuy2GrYBy7GfL8NyoKpaR/TEBTiHF1
eY5zMvpN6QGxNe6wh/fA3VpOTeMTrTdShsYb8NYMaOyuSUdV278XJEDQcf2BEY2620onlzRRjcYU
UUkbyNllOe/BP6NSxT1s4LIWPI9oSxuOJ+kIrRs1tYRZjuFkYwJOYRSAShgaJBAHyp6Gc1icUhuH
Bf39yCPQ0ySUC53sXqX2hxpHnkrEvksmla6e0Y1dSbzH+6YsKoneZK4Alh3aDXWgtcdm3Zq+tOTd
Eb0C7cx0EIwBdZihNUpKdESjJOkADSC2XbQKdLCBIkIDec1s/xeOXSlboQ1UpM2+afYbdE40/3j1
uWfqj5TiZcsMXMFvB6JWUXhjWCrcGXezDdczWjjNts3VKUPy4NgQVDfjPaJLPBrg4+jH8mkN8xIq
yk97CKbfzQEGGu+/6eGHsFo4Pc7wfC4K05AQPfJAUXnvpxt4wDClvYGxvOikLlzppxBYhyMJKbhZ
alXHFJd83GvMTBihyHxmUXNpVINz48c8Rre8OIdPAfQRtVm8HpUYwi1kSKf9y+yyD9N4ltnIVtQj
6LxTHZ9mn0vnXZQTfJwuUAeJHMWEFadPfUsiHXlY2YCtpiY86+zk64fznkmN39CAbXzH4P7uI4+R
w8FgsAfQKDlj5PeR83I/klfjuCTDXvsxKnCfcRPOeJ1Q0qn9M+j9Hk4aamJd3TK11QR8GKBJTCI4
n2xfRiTwBU2hsmexjfxoJps2t6i1dHxGYZ8+O4MdbCfqkPNfkGoVdzBvUHosBzJPBFrXYxeSztkO
JYExwo5WFxm37dTWiPfurAzyOtmXzd5tdGRUyCMsm8Wb3rsvEnzU/xOsFc6CR1NispQ30wN6w+Ng
HrtCFnngZsotZA8rqE8HFxQkiDTmBfXEhcKKxr1tZqdyGMOYZQYR23dinlddhpIdOF01D1UbheEd
7ADztsWRSxNsNad9C365hZxWx+G9++SYfrL6yM0DYAVpGCfp6szQOuHvId9x1//sKVLzpXwKTiq8
7g39jFSIa7quE03/uEAr4fMK0mtRknbgttDLFmhdeFUGXCZEi+BsWSAZx2gAC4Uci2miVEuO1bjS
IrzPIVZpIDEyRRn6bOlykVhbCwrNUwd0nFLI9NTQeXGM0YS01LwYcEIHwRg7V7g6GCbUC6YQTSDT
bOXnEoyLQMl4Ud0Q7QltEqZAqizP13c2l9TpQBVOl5O/M9OlwBz4SUwtD0ZOLb6bpru4hP9otOG7
g9va5WYSOPsA7rCZ6B1PlfCRbSyvEgto6GVD8q64SPfA6ZMVOi1fh6Mjkw5Rm6cfptz+byabRhWN
WAZ9pxEyo7sO6BPr84GWdK5oPrLF5UTW2K88Fv+2GeS/jKf2o3K1tkTQbO88TQv6LMj2RFr3u5Of
1O12JZh7jotTy6Y7yq7RIspqWlRCKtsGr5T79oSsBOGZFfxW1vahJoMtYDNmfXmBx4QyOZH5VnH0
75cZ5pDaTh1AooRkEgETC5WVvsEfFKOeqDyT88kQtXZ+G/IjrqQBUXqim12IuUYPPvtOEbIoF0lX
3elYWMwZbC1j1IvUBnHgG5abaLR3Vr+TxXLxHdv1I69lnQiPPGefIe59m9w5Mc0NVmHznvpUY+iI
GuqA4MlsdCv325rZ3Lr+7RSy1KZGGUvXHMOpci+6ZuKItJl9OzA6wU+SrcaxFX41mUcgYXnD/R3d
36VoBCwBnH8gCUvGkgnS6fKxuciNQ+vcMI5NnXG3gN2QtdXCVZK8CfUs7mK3edBqFSvHZqRsW0oo
zz/0lrmRCZiRjotc2Ug7EV4Jd2t5aEZvfGB/shP8Uol3hrc1E4pGSKSoEUqzVNvSaWVf9A8TAFtm
eqgUzCrnj/ieWFHLXKAcqvD3cmALdOM0D/b3hwMt6+smQsDA54AgHPDC6if6Hh8X5i4G9Nm2I9Qg
oUQ0tjuykzJYPMH1tYphSvoWHkl5zEgpLfrJFWL7VTgWebSrl28QBFQ9fg10ZKgHSctMB56yrz4M
46lcfgnxr6Atb4FHsesD2VbK39LUr+N/EQBiKp86H6LKnBaIs/QSMS8dxvrVSocZrT+UQ8k6BYG0
OCN9yry295jjIIqc5GVx75SQOHIAvmuVHwUET5uPGTb5R6n+cgaq4N2L22oWy28xUnJQ6I7HZy/Q
dW2/Ip5Iq/ac3QrPFYXrNRvAnURNVLV5n5PoEBUnHmCTwfCywzk25rpvKLfZYTRoBHYvTe0dw7xk
/Mt8gAKycXD/YExHxxlXAALn+lSfnU+Qd0TI9jcEEgoGkWvWKb2ackkijHBceC4/80sqcNslRhTk
grO0W7t0ufcPrCEjEDfI+oF/SIxRUn/aj57x2lflJdGju4uXvrdTHWkVrEy/9uQbcck/DkT29nLF
g9N2x2Ql2M6/M2VVyUEPe494xwZDft1lI1gayzX4xIlJnr8w/Amx4/3Z3000jVVyv2tknmTFwER1
kkFCGt0lvqAmtcu5cxntHznSgnkSLRKQDMiZdtrtwsS135R2VM2G5DgetMlJRN3pIdo4jtmr3NPc
i7lVAR6uMTgPP0hA3k6RqDc3HdA5oXLCUkrDn3iszoYhGnBUaL8CIMF9HCHw2kQ1tnINkL1DCZfP
U4bKGdD6NcJ6okMqUeZKFgdH0Ukd+eSwmaQSPMuPSU6VeVGx1bk7PTe4Vy+Sun63EZdRgqMq4OOJ
VHawc1HJFQXsMkBJHa3rBTv2JEdi89g8Xtb4/ugR/+jD9io17z0nu1K1m4WUhQhDulxMJQofafSK
2jlX5hsCsUam0JBQHHhXJYE4Ox4p+7U0WXLPCtdm7pQkRSuiPSGg8tyvLbafL3Ilm3UrojNzi9e5
kc0JpZJvLnCptUhqiHCQF0n/8GrZEEA0OCgvkiLcqgLvl/m2pZWf0q+RBhgoQtrb9TF0tFKVpWBO
EifDbSddKD1bzV9TmfIQlg+Np0wl8pvWkko3ym5lwC9ZJz821ohCs30ZR3kHhk5F5h9gwFNdea4+
6bkY3mgxvzpJlQ2YIC8KfFWHmg+Z0LDHXEwCaGE9cTIy0g9UoIhZ3YIKHbwq4eoidv4/o+dV6+Ae
j36OimgD6RA9wc5TaObwAp76N4zTvhiRz551oejJQZXck1/Vq2DdNltUtoq8+ALvgLhKSSV70qX3
C8mjKlDqQQUz+aE639d0xbup67YTPkf7/1i9zkduIIas0UAs06m804SRWFOubDHxJlAeaa06kfli
HQKs0eI34WG5wa9Lf8YnVZ7BZXNyKgGy20xpsW4l9z+ptwMc0MQG5WuOsGIdqlzQNn4wPuqODf7O
nyhZZuMGYlOBvLs/nPQYdoInhX12iJxOGJrQjOv5L+HVcpfI7A262zXlpdNxrD9SWFUExTvmoDxf
fRYSzqBs6Squj91LXFDfvR5VQvtAmEYhey3pRrwhxapiZFZDeVEqVb47CrkEX2jeETS0OcQ4N0CB
K2VbgFjz3YO4M6SvCdRrMxhU4lGq/JqL5oHJV9xz+sFlcWOFBmwu7IsEJEYy6Z0IBpb+2qR8UPyT
hXBv6co1+WQuz6f5xDHGNF5L47CBGDNfo5GIYMaWCAJYOsRO46xn6qwo9XblNqismIAuReCcdiRi
ngs00FGiFxJJKbldA0SDBU+RsLMfNBsgOW7iV5pJ6tJ/2g+o7rHNfvlCCQafM6lqvmnGIlNqdfdM
lZ1wFt0YigMRNwqwrLZAAP/IElCZy14lgNZZgGI+Rvs4I+ytZEA8BNnmzBlJYZdvUKM0N0UpC7MC
ErqGTEEjk3nUz+IYiVZ6rwvPbuhxFJYs3x7v+fP6qNzdvoVAGqSvJ2I7OQunSIRbvtBBBY0FqS6r
6+0ndOVeNCLI+9S5fsJqf/0WftbNI3UUEBC/AnJCZWuCJllMnQWrYJwBlzzGOhn+DLZi1Ai5BjXI
6MVKTs2FRuOBkrNb/YkE6X7c+5q/El6HZQqEJX+nxDEjACZGBp4CHhG05spMwFKpuZlm/qQill8v
PzrxSbAuBkYRC+N3WFrjk9A6/X2+sdQzzOp6U2zYI2VSz5zIs/xF2oVROfn/bG9oXJJ7sOjjGJEf
KcUZB4XrYj2phcG8//X/uHuaFuHG0S9LR/ttlqoWZGytWxLtOvSPcVIN5moViS18RK2neQMSlgi5
QjifaX1TZmbICxQ4SPZ95Eou5bpVbc1u6ezT/UvmbQm8ATRKEWkEGe4jLsgx0CSiaSTaaksXo9+7
Tzb19Mx55TYre2VT8ipYV2pj4TuhRjmP8o2m6EWAabeHYOrrxyl5NDMQcYyoG4ynW8UW4Y1jXCAi
KBa4RH6b6g2YzDiukgiJRvYbEVmmhNGm1+fb0hkwilQ4A8NvvNZFyEJ//SW/YRfsU43iiLEAXVg/
QT8Aqhpv+i3v9EpOqbgy2fZBhIsh/qf6YbuUXl1LJ+L51gly9ywPnomEXA2QdAoIAALqtgMj8mJZ
erlh01Use2BUqfFq13oB14AAQFND7mHvofikFUef85pIt9h8juFqMFSircX6sT3NWkIFoxzzS3p/
U7FtF23n+pzaWQZD7aNychEJDT04+JwxNxaTW91t+x0lZuSd3Pdl/rej+UbRT3QWiQNKikA3bl4U
Ke2NooBh3Hv5ho3by399xzU20+ng95cb5P+Nce8YIPD+ScZ//ztLkmiCJajdamg+EWUnJ5RLIj9c
++y5WVvMMpY3naDjCmREuWqlgrzEIB/UqmvUoX10x14W1Z2r4WaQ5oP4oOwgky6p4aLSopMQKElM
fArHnLBmaRRWGANW96vMpD8wsuouUDB/vNX47I7Hc8evyw2EFfpvrZqwnIqrFPLSMPcSXwunp1xs
2WFvdv/4ohan01CZJ8/mOmfJsHjSjlLdsKSFH6QzttJLMjKqnbsaJRkd9BjR1o8BKhj/Q2c4YfDn
IFcy8QVgqCb7CKvu/vs7wrpGs5k5uwrtLulEd3XJpxIDe7IEPD78QXj5HoFXVgl2UGK84xOyjhSs
OJxD/bcm91D0XyGtmOXo+DCih9GkOzhi3ugMLQXxGt3GaE9pjPEJQ8XEBxpFUwgwroD7mFELbRxZ
m6ZSxgbETFWwV1Ub8H7lUK7foGsC9c4lChEKk98cAnctWTnNjQ85S7H9FqU5mMwNkf8WU2T3hdlQ
CvvxKq9P0cCRwB1ydZN0p5/3kKkvrdNtyZLxBLB5j9gGRAUfoSP8cP8zRnLZ9i2hBk7h/6KhsOy4
/ACBKJZvYvKV8w+/6IbZTaSaUBzgUoJIbybZ6G083Tj4gla08v7US8TrOUIOnfxfeG5H4CuPMoPC
NIQ7zoOY+Cdvc1/0gY/0+Xg7dHsWl9BHstszBXu4Unq1PRDgwG9z604/NXt6eo7R7kAii4V6ynuU
oEVauwv4NC6uJjTZvbFDHojn9yHDGaiC0+NDehH558qICw7Hrf08yPiKLlEk/ziyzLiRPSuoY6Yy
o2vkGHl+88v5uFImX2Z41CwdNI3ogRa3wyS67NA6fojfytB9C6sLmkRJ2NrdwO61sJZAEqJzcF2X
4RHvpqHLCVuqpVpBBanojygIx98SLK1MomyC3X8H2Bg1v1Sv8BIrK2YfA7TGzMXlHL3qcy4aia0D
CyVUzhBot1x2sFFM0mv5rcYg4Skq5cK5Af9E8aTUftgr52xr/5uILc7YzggsijM/OGADVpINJaVQ
tuhhhY8D/YDX5Gdqxe3IufqYtWmGlzXk4cerqEP/JpehFQ6mEZby4GpvtqQE+DVl4WjSx023qyTy
ZWz8/5xSd8SfkLrq9xOx4QTA1miAHNfqdQeaJ+ij9hmfVQ6NCY1DY9xlqknnAMxl/TqTFS/pSpVa
s3QoU3zq2jAJsrZY5WmsiBIoERMdyoxODskBPZSpfx6ydWSj0ZrY8wOE9Nzmk4TxR92zKvezVoLr
3X5hwD5ox/gkq/jL0X9tklIytOigolPo6unv9vcDZsI5r3j07MLTcSRxIvxZks3sEadhRat3Qbbc
j/GHOJs8+nkL5JWO/w5tsUGjvfjb0gv/oLnV+3BaOmwMbnQRsT4fGW3fA1tOOvLwDL6Pr5K7Hs0i
p6XTeZsbMKxzERU7NETHZsLRIc+FdUxcU5sk1RcaNv7BhsFTrIHYCcd5W/wBkFPWQrBR5rN4oQma
bvt/vXSzpLv91qb7OX++8EjnkYXjsUU7Nkpv9doUsds6vql14AyJUlG3j5we0qnp1BueSlfcHySF
ShOh6uKpeJbgAz2pXPaQw0GjmqpgpADP7iGk418vuh0ZN3O8P1LwUxKwIOHKy9dHgTQFTa71D5WA
vNQmG7USii7zZieecgMbqj914mtn//mDLk8ulL9tfJUcK+1ctTde6CSQ3Fc5FrDOBvO7W/ukoJQz
BAZngZRfsdw5FDqcU2m7DeTkZs5+kpJqyRLx4/vJegCgKagvo4/a1MUyCoAlogwM9fl6ObIW45AH
Z6UG0PR73J3oFcydmgGM0URGF12R5pyW95D7N4ml8YYqzs9QS0/3VjStVo2A3kRMgrmV5syiL06u
wklxVOmuOuKMK/oSRRGSfmj4wKW7Lc3a10NmXsiebjyps4BAFiO79+tydfNGFw7h35XEBobY6nQd
+CLBHYlCNVvIhEfHT21AXe3yNPL3elaak+YC+IuKKZTxIAhMgeyTGn4KNzYi7NDysGGNJP40aT8U
6XUuKKgwuHNwBDiodH5qE9BeVTYBZVvfzAtQ/bimLWawDwZR9iepT/ijZqUZak0PShFJbPJP9LZh
Du+nvGPUbS46UJWmoueYG1WCD86lw0KZw0VTDtm2HgLzIJ1b+9rFKjVLRkMVfOma0ye0RyDuSDwk
todeeXeI9HAvTHgz5gNiVHMwQRIvjXt1bKvJDo7z0x8me/ZXW7EQkKpYdJo6K8bWcNHQlRyUq/FY
7UjEAhb6mFONWo2os24NoOcR5HL7nQP9rGCLNe1SLYP4PjVJRy0GhnnyCULorwihPQ5Pkvbd8Cdg
JEU1KwMPB/+gmSAYUc7Ub/vmnIqsnGBTikiIQ/6T4nGVJXFoOwKGJG/Tqi05DBTNZQfA4OWrbdu1
ePANhDdgCRysrM0OcQ2QtqU7OeaHzzcen2s2s8+PdvjCeql4Rl7qI293XkrdeLOg/Q0KjjtmBLOt
/kXyTHw23R6mTkYUbn+sPmypq4pLdy7btL8bVDaF7Ymun2ihp2XOA6EOIEA3tuc6maqo+xttV9K8
qj2wISqClTehG1y1fuE9vA3Rb5hKBBAg7HC1YPnB8Uh8YYaCPPUInxJjvrot3wMP6tWZXg20tB3Z
8+Lndc9cDH1SzJtY6J+IFMxD1/Ver2GlcOZhls2ZzEsXxdjb6bflv4nXPtYEhU89B88FGUeLi+vJ
B7Afe5HSDCgGyZwC5xOLkKVIkvoP4HpWWzotQnDfOQ76Ly98MUOk2SRBwFeOSWoWJ5mdneCohp1I
HuEep3wC7O90aiuoUfk4gt99TSlAb7Y4Mx//+3qQMQzMBJZ32ebUSJkzzyjvuze0ZgQ5udmfw1fD
2xu++ZGSRFIYs6VhqlFakJ9D6KSWw2fvr/bfXq9fx5b0sqxBtLcYdW1pjCFjaDthVk1OQDUVjlB7
pWShv1YZXM2pZitY0fDU2tPLo44rZ2XJG4harzeYcqtEZP/J8iSA3zTuuv/K12PcKX73DREhd7k8
/mUY76ML2RvsDschpVRqc15dBHuwhpep9rdaELhM7vPS6h7QDNPY0+fWTSTDwRQ6+ns8QIPwbmyg
+8mVizPNZ6p+RLNVpu46uOba7v7rNFkgbxKGBy0ENQRzbzarMd9vCi9u69HSaHM5kbzh8IdXtUcT
VCjTJBFpfT3cZtRsrp/jW24BzY3qReeccZviJHVeAD/YZVNE3ifKVvMaDVyna0pmjPKH5gyb3Bpe
Efa0w4nCC3jkcSBvajbzGtbvvmv6UuxxUs7YsJwr/esHl12mUFKmxUNH+MvfDVO7XFwu5/YifsNA
ss4A6SYRBBP7V5ylhQzuBZvjLFHdrlN7c7LBy0d8ogZT3R1FeOewVctcpae6L4Iv3F8RS6Hsyfp3
xF4yWMAegUCsmquDVj8j6i8of7KNzV2ljQQqA1iZf6zdG5/23cZEUiIws0uUrhzrotpP85jpPBQr
jo2fHynZmvy0QeHFYaD2NadzYBu5lqhx33ldm29zFyAm5lfnPdyHFvgF9DFaPOFm/42zKleD42Xi
yCrMhgDrFP2rKZwNCF6+5NL+YSKYKpY4jdDuQjxJX45vZU/k74TNxbDlzjR/PjiBXQDjNB8+hEm5
vDv/zFQHnbup5fIlQYYACeS9Ap4EOob4JNDXaGe5urEduN7aOQRh4yhfjsoGb9WEnFaaq34Q6NoT
SkaJJphkvgBTPp/lLDXc4gSki/v6BToPN/dyTfeEo8/gJwa21xueq59SXD8F9E8mVUfKqR1+R1Xt
5flHKdaeqUb5gzj1I2RUZx2CKpmSH5YuXp8yjq5v3vdW2n2h3/rwU9MDc2+ZRr7Nl3K5qXOuN2zM
WGlcX3xeZOoziJXCSBavpmkcZ4wB7QA1w2l1l1cuF/FvwWXw/5rr+qyr7G77tL0f5ymzrrbI3mOl
gTP41neaXlhT0Ad7s/0n77Yv8GeFFKdew3gTBv1D6yl1H8u53/oE/fJDYfw10Ytaho4eLcWFCqno
dHA29chO3Uj4gQbtNhcKVEJTdfhK4L8r3Yj9qkoyqW5QYQwAKtw/VBtFNGMl4SPTRAFYWc8cWFeD
CWyfpnq9JMMg9imn0NPLiJL8ED/Elw86cps1TB8M/TM4GIIESD+m6aGmW/JsqLAlyRldDVhdcwPU
BPRWKsPiPAD9rSgsg2mqa64xRi0xxpY8i0cTa+JvNLyVbmDyMwinFu3JdXQa1aNOwdwGx/4y/CLD
Qt7ZREqAkdU6OZEUEpLRRU95gyM6FDTfVtIt1UyGKP8CbOHNUtwLc50Uv8espepBxIA+gw8sMWOp
uH1jjzCVpJ64RCMzsVysmahnCR0Imr1PXKi/2ilQlTUfQqEEGgzuPbSaFpCa8t0rqqW+75fdR0vz
B9zGdYG31ZnP2yPrC4669H46OuvM4EyI/wZYvaLXXB/SF8nLTxd+eSeQJ9d4ovuUUrXG6h8H4Axw
Rm3zkdPjG5jIjhFdwSzxQwkr2Aff7IdP+neTwVghfgkMbCrX8GVg4c1XW4VonkJ9tEEcMSrHHXJ1
ypEqpd+EMOiHAmNvpUWmpkiGTk0JXJFpNwKSbVNm+/9F++M4tX/m9X2IAxbS9DwmAzrOh9utdKuN
JU1lZr1KjPQ7PvUEI1r/jw2Ijyhx4CUn/SFyTfN5z0WBN4dKvvklq0l85+tjqw2Vj8CKfZywN7rM
dkIUalSFKb95SfyfLHqHtKAnXkktwzT9oA7BznjrSCKZA8uXJN013GtoxZkoC85w4XHvx/Nq6lPZ
CsiyVKjnxH/VVWg6bp2PizGPqPizxPAj+sfX5F5ZE+r/8KmfzggMoUkDOXDCC3LUcEK7h3nxGzzA
N6exD7dwbOGBAFPjRIzao4pXvZoW5gDUS3QRHarjYvKym1v+CPeb2VPsReKL7R/1v70ZlgHqKK6B
2YQXRz++orVYpRoZpOjJidUwLecI0CkAEx2zQNp34RpB/geA0VqUAVJDpo7XEZvoViF+s5vDBel4
m1jV1CZZJ2fI6mzNOvRCb50r6g3NK9ZflVvHqxnZKWxfDhJhCaujPuh8j5C0GhFUveA03Ckr+ni9
XvRJirqEVI6InRUXmknWkzId6JBqKaHDe+yAJ/fSKCLV0TY3XVSlPCC9t5bGZXaQaGKFTls7+kzI
SI1jw/RgjrSkb+iIMH/ulEssru/g8MRvW83ZpFJ0QRQ4STzp5cE2OkjKP4khITNWxnft+WdDiqjK
ImQX3+tV0Y5BKDdyM2S6PAzNbZhJTCvD/ihmjyu64Q037JKmtrNa1pTQl+VE2SAV20/FzNIedB85
KSVaVp/kHA1n2EIzGAhAlG5xeZlDZTk86oxJDdfWtHfcWptt1z1vgKmLweOGKgZRU9f6j3UODZlh
QmTfjkkrWkKEyV1r27cNn1VFRF3UUzSMYfHwDAyWPAWVFtjWAqa5Bs45EJYd9JcCnAzFhb9mVb7W
Bv1XS72CQHG41+M2bRxAAS2AHdcfbjivSy3nFv5/aDIfvU+0alWlH4S/07w/Y5lNpTsKKIpsIhPG
yTVuZ/bl+1tr9beWgKb8QmqrIuWn5UWruOfSI0RM+0ymDdmGovbx59JioZHikYJZv6nPcaqxejwP
WhvN8ryoV+uh9g0xft4q2tquSTn/fNbNDUFoksmgh9POpZaRqlXIJTD6qQkSxPy1eG6akJ7fSq5r
3Fb69NTZKp9TWvoTUCyq752XaFioP9Tc08REV3S1W20ucm7ffJKjiHUeTkeoO34lTnQi1YtZz1gO
e8u9v2NBI7y10UfQZVyK0L1WIo3Gfr9UX4tHrOzj9qcgPQcwc/XoJCkaOZPSV78vMXFqWf6O63XO
sXZQhomPlOelZ/7anhYuzKGD5H9tmdUEqty9vghsAnUjMe3Qrc8+PTGuaDFCq3MyyIWbq5vvRmcZ
Hx6EG7E/D8xNH3/PyE2fqipQOJVZ7GX1uSWVhOIZuflxItnHy6KHQSBmUajmzbB9SfYyfO9ollXR
n6fNvBoBAGkW+WQBwJD3o8Kp6Vq1pKWfYhOSYdXqY3mAZZDUlyokB7aesTlP1F3mYSgAXLmMjMuf
RhQaAp0UxjW51UMQl5OEPteLyzG8swpnJgfsbHsrQpn7RwVThGvLCVo/7H1ZuJJnzLuSKHh5Knu7
FKgivLBagiYnwNxhBm9XdyM0VxhmUFhHummZeDpnFrnuJsP/m+lE7jgMp62x/fg39orkUcTT2LPE
+0SaRKzw71xYR60YfS3lEpPtaywhxqxb23iD3lV7nV0oMorFexyplk3U6fGsLuxa5C3RgK04meCL
VC8Auwg32WCm4FMCq97cq27wg+6dQ8pbEIY2WinuJ7OFkbb26bRPeDjGBQO3LR1lj1h4CPg3Ftsh
Pr0hpuuwYVnThTPT2fiMtVjWdeMpO7oqq033MxB1379rP+KeeVMRop7BDwwZ13cHcPGMxTSwGYPu
yH7MY82tikOB8c71H9w9WPGonaxQBy7xxzXK1HqSdb1hipbk68c7ERayuj+7oxOc6BRtcjarG2HD
12jYYoqbnA8+sznUMPUeDOM84SqW4CubT3sN6Mcv1FyHX6x01mYiYzjIeh1xyPOIQ9F4Tn9tYCbF
dJHPaEA7O8mMYXR5R+qD6dZfDJ7hQienlsAb9EG2CjgyC87gLe4qr1RuU/bR1foAQia4gTXpG9uG
yNoroagCxnYKlJQGtyD5luik/f318SJc02f3Gvlr5u0hOrZrPAIduhQL+Ml+OkDUXy2wBC7ug/gO
u9r6vTAON45V9fvDXkLiqq6w9MBC5Eg0pF3uTBXt1muDp63fEnXw5bh+jQFmlNsbIZ4i/P1uOKbi
clEeZMR5C3/JmJdswbuHotq+uT5QJ6tjHW8MhWyzgdyZ9i+NrjvZsguDLbKaSeb783FISfbxJ8nR
yCeG0FGYl2XIYfnhhOItblUC/u1CF7Udkt35scpsmayrIPDUP/8GFT/WnKxA5ACu+0wqE5QJV10O
XIo8bppDJlkyIgm/gFHGsA0XnExNzK4k/0Pf1c9RInDXwFGRtQhTKRpkvCwnGIVlYUs6iXPa2lRd
+XiiGXUAGFbYJvX1RDBzpS146zQk1aK7UP1Zis1LZfmgn0SjN5QS8l9f86QUs2d5lva2bqJJiyvD
UVdoqjgvIkiAjZsWl2KhaYTWG7934PNGtQJMNIClkr1c0sLK/Y3HB8fPRc8Eq1G3uFPqS/2GKl/7
/elTPn8l9AYwu9SMXclSbEDpf0GLMVfb96ABf09yUym2Tghk6sirzXdRZSmYtisMZm5B3Z1nyLqo
reJqL4CQX+5WjI5zT643cZLWZJZAeUrd3Kp2aP+RlFxRxyPyJDf29MsMnUqPERZm7wOJz8+7A+ql
e9Jz4YL+SJxbLJkg3copnfbP70isEQLD5UQSqwbf+XPTBuk0aJz2ZN5weDJVOTbJz9wYN7EoZfZZ
I0OYluauONs3A1d76CaKobQWAsPWHQADMIdput/gOxlAz3FDgdkASnxUFnV1UeeaE3hgiIFkz0c6
84DJO9222+oFaHA90Oi5qpftN7aZpSbe0OFjzgbGMq4ssQZ6SrE/RezprRbyVHN0P6PSJvRueYVC
EMSusgDve8uxbINZhJ9/cWq8Re0L85HvhN9g/zDeXMQpeHLCugYe1ekHdaPUVrb/KDGwx2P9plmB
pJpJFG5LY/0K4EVaUkdo55b/3Rjgm+1QY5DHWCeuRJqbmXyDxivPW9nGVGZjkkzKCeuu1kOpwUQQ
o9L/vfNSp/pNjdb6augqIcpHy8RVWoE0uWC+xcSCpS2p7eWqILVIhPxzqDQ4zZ19O0vncGDd1ZQZ
my90fb1ekGt0lhBfocaXFTuHOQ0VkuBZCFEw1EwvIzw098xXvsSXfKr+FbffaRTjDsKD170g4iyG
ezgFHK4Y5FSgUqA1gBt07l7wCRlfEi95bokvj2pTIVJfzZmAytQqnQoxhawfniViEO8e9RKToHWF
pzRPTf7SK1Xe0xWqL5lQpetANidrETKMNGfpLGPHvaaurSoPMhXndhvs0sDPbgBLmxf/4ymNrfAx
pkBZ8rlm6QtexXE8mqnvN7mCbEJFc6ewFWXyyHMeH8w9dV3yNx+zCR5cx3SRwitXgJ0zGOkPSKK+
Olfja+1aZyXXNBk68Lxcle0W7XJkMuMkug3mD1eVPkA2KkcXcee+Dg6RIYNFGHvYaSG9JyiklxrU
x3qn14pTLB7iEomtGJtS2HymuHDJSXRYgkUI0HTwtWaHgaPz7tNbTij2OA47ziroiCvqw2MD2Ocs
JJ0K+E+vASJZAfM0VkS8lBulL+hznUZm5GofdT8nKU6gUFcmyW6vrpTydGbEs1WezXlQyCfTV1Nz
eMR6SybhqAeC1u+6n6ac1Vll24KYULnvvzafVewDbrMvTSLFXb+LrDzCyPNtaWbDb7gXQM/HQJ7j
diqrOonoOEmajgCuPo2loZzLRd5nMS+SSaRBtJqBs5CQYTszRxUElLlS916jYqIeybpk5X58xYpP
4m5e8dXe3I703RNwU6jggn4hIFcg2g59p66DmAG5Zdijcoh4Q7nCkKR5C/73e2cC+eMNCWpsliHS
uzECdTW5ZaZe8w1JUxQdWSxZCnwVjzgh3WQobUjaSxOMEhJjl8dl0WmqivQu9szATQYTWlXf9qpo
kj7ZGhulgORfvSb0RCRA3eFHpyTIecgzA5nkeGVrrwl+8l+tJr4kPBvcqCrHTvZL/sCHmbGyPyiJ
8f7Tgh8W5oPUWh+04Bw2RC3kA9xZe0/NDMu/dmmSFy5sFOgD6TORyAivtv3H3YbpASTJcHBV1R8D
aVWEGvicrbDt1djhi/ceWiDnfpd+dtZy/NLvJAAAHBRR2+DL1gMQSzTdG0LNqejgY2JLmD/87DN1
AQZA6RYI3VfWAelKLc+w6aEESBFzdBkFIwjdm8fVy05MUP0Eiw+/40EM3j9S4PUfwoKQnUnR6CWx
UWAtdTmfJF02UqpAGr5ehLc5wN0dGA9qiDi66SW0JUbnvg3TeeVSI4TJL0xdOC4d6MDLoWZDn3SY
eVA+q+iGUHK0YZlRkhfh+z2s+NexoyEB4iarUJ02BwObtblyqxnDEP31ZkMuEy4l9tIh9koyaDXX
70lE1pbwj5gl/6NoPQc6DId6tqEqCYg3SPxX7heP2OWfaxStPsXM4+dlTNZbK1VepGgg+lLQF8Ui
zqvamoNAIN58RhieDziDFXQXFdfjuFw1T+LYasf+1hJdKGr6XgWZbfJMIij7wuHHdys801TItWuy
uCikc2NOmtbdUWswV0/qtg+5hIpupM3o6vn74XVRsn2rlb4AgdQPJ2H8ZHcNZR/vT5ByeW/6B6/m
OadBhaKvos0S7FtZcBe5Evv01K+n4tLAZpIOa0uEZYD3HvEc9N1ajKdcq23z8U4Kx1/I0unrCPFI
oWGi4GX0PTB2rdV+8vPsP03kJirPapdmPUV97TRXylkIjXnTGkhC/TehivkpMd/XX+S9iu5XTnM3
uB0tVJ4oSDBXQu8xLzNUeYiTo7VGJ2sohwhr6+IjO8yo5FTjCwxLaM71POv3rv+TMQGKMqfmBoFo
WAECODsTwVtrpTM57mZwdCnwMkMRIOrQQhMwMJo7hhhORsXagSivYVa/nRG5iGZATiuCxzyY/qy0
RWCDvSIopFsH87i3Gl+9hBoASEtuPJs7K//azGOkDyXWgU84IrdtJCGXmPJmXODGQ91Nzbcco2Fh
+OFPnQIfLx8COR2knH9lfOVsLElXEMJtNlee1BrO9x/Be5Ny1d9IsJPVvKCOUk9ex2lEHBafgNCf
BN8qgAS/y/DvlqMDyefB91uYEWT+3V74ewFs5BJp4IG0hW9ILX2/k5JBp3g8iYZgT/014m1uZ/ct
y+p4LHeube/jQXiwB0sutfw3QWGlKkCdR4A3xG3bmfODO+VdFXB99CMbuavomFEOMpP/tODCDFqX
DKw0wu6HgCOWII0KWOCFF1JdDSrRcPQMachCp4uLn0XdCkOCeK5ijdF6kNJBFeUXuQaTMXgkYcCU
lNDkps6d/QTeRWbcK/brk/9UMKtmcm5r6bQD4ca0oFiK3zKwflVT3bz3iIBJHCXv3ViwNbt6ALXW
6/Ghu6bXXWR52WZ0khVmyN/jPyoR97B8m9MLj4DOxA7WT3zRNferSLEOjwZZMs50sJrFLCP1EJAh
/PQ+6C7s3L+nkvaY8IkVd98/72EL5x3KrER40Nsf19nJKr5QjVwyzll7tKPNk7sxgon1nnOmx6pS
tIgljdcFzVfpwAwmZ13P038yO8qC+E9YChrt65Zhh6U6biipqVIPdzo777bqjBUgOKGN25CrFrmB
qLod1z08WB53ZY4qiehejqTA+rR8f5e9qEJlZbzOnRKCmzVL5eS0L2Q1fE+u/hwUFF+EPqOcJC5c
sZP0FGwBdpFG3zNUHjdx3Q5Rp5hjBvVLL0YtDYhICt2k8TaOPbpvUauYAdtVBhTkUnHRGqlGkpig
cSrnURrahWVRvD83VcxCYQ4obtevCL66u8okoGPWCrcJWWn4QmqUeOy0yG/fWZDatL2kpZuG1RIo
vAVlNhchue6GyPbxjYughEn9K/UArQXtze5K3l9WllDhLebSCa0b2OJM9MwFFPg0GKSOg0zuQm+z
RmJmxnE03kWvyqxU8AkjrZju/kHXn8++A2O42QpadW6dUsVTrhTtJLfIvbGwl9H/rtmE2jFeHuuB
tW3RnEyTgL6i9qiNPUp1LsYIYZfOw8Fa+AJ3ZZzfmYpDXPcT42wrMKYznvpin+sUdrX+zKGeGLWD
X/N62BJO1KHPGFB1uKjZIlm3utwKpdeBW/uKZ0xDY2Hq3uireWbiMVUA0/ZYv7klzFrjp4GN/KQN
fjS3sHsuD7pWaqp/xf9hvIrIHACLlkxNC8wJUr8VuKWYTFM7dI5AZ8iqKdmpCNDNPL4ZeJd+1pbH
CE0AMfDFidMMT/6lusncNAgAuJDHMeXo7mN5qnDlP8vUYpezqOW00lkZuipwgVDxfUcDnkpRUuUX
17+pPo4TfG7tgaYa/SnQpJEdGQV/VSgdTW+Y1qY5njxX24hK0BoSc2VwaooxVvZBBo51k9pDOH9k
/dqi42Tzow2Zbe53RmQKPMgfyQJWbudb61oXe0GAOwuw5U/Ln9Yo5vIwCnyVIYlRBeupYRRt0bYV
vp0KTsp0JzSWSb/PrzAavwVgAtN+6jSmi1S//rBVooc/V40Mwyxn71FpYeEtcgZhJCibAiukF5xZ
/1ehiNJY/vCm8w8A0Nqv6Q7P3wQteKxIeE5fJLAbWKN8rBpCcqtk4nV7QWNW70hgw46cVtx9j9Rj
lBZk+2wtM2Q/m4aBKlHVt3YzFg0jyvvXZ3BGD0cDOHSgTcTZksD7ZO5/scAcbVvPU8030p6pEeze
jAX2ArMdmbX1hdRWkoqdWL4oPy4WD1qrrmBx9gGeDkHe9PdfgmvAKEcVkyaXudU6tcIfW9qbTM6e
SmKRMd/xN9Xy87x57B5Y/82S57WGv/K2h+QagA3+Ig7dw2+35JFfrms9UHEHGyVE6+rAHTPC/11j
qUx3STlx/uVEHNqbsrgWiaJgXsru9b1Lhz9h/vHGbO4cMeLAsC+F0Ty1428mBgIVP85R81pQMo7n
Op74elQstoqsrLVY04MIolmxzqqo89Od0nHfUeoKm/OZCL0K4ZpZSJT1vuWp+F4KqReRQ2ynUDs9
Z0sosCQhdmH9DEhydOwaXZAXQ9Ykyu4lVOBiWQ5s5hnVS+AMIWgTVOAoSV+TiO6L8C1JNBB0PLAg
Q54jYbseTeHcUgGeljehqW+FekTduWAcuJv7ufcr0cRI1kBkmb59WdhfmoB64LWIp+PemtwI1wjr
EtVQriO3v41g3BOW6WPaKanro2EmyYDNsFt7y3wJlm/ALzcMelmHJvO2AKBuw+OzNmXvN1vi+oLj
tfwGvDjc3Qs5WLm6MFHjAjhZxc87+QG6zBk5n0DNmV9MZsuXxepjPQ46ucu7HH5Ve1BbebvJouUh
RTjjj1uG9Que7WYwU+QSY0N9aLOv82dvd/Cymq1L20SCm6ZH7x0EYSRYiKdCzijYVp0cRf16B+EO
e+b4bE9BFdtURgmNRkLIRDcFr44ErFL7vKLETBzYBSQ14oCxc+SD2AYlurw5/6olyuCl4Kz08gi0
jU7hswGBL12ce48jzkI4jGKRA12HU7lwps8R2kn6CYeNJaQxM9Cb/jFyVvcf9VkBJ9Pc1uG3KTLE
vsfkYudx8JJiLPS1uUyi5Oousf0rt3m+k3pqutoDbqg8xy6FK8//p8YQAGgJb4leXf5tUxp/7OI4
UT/XEAJlW7CP00N32uELOFElemZusx28aLL2FZeMvsjLKJEKzuw3jFwQnlBTi4e+k6vseaAjymsx
FnHvpZmvL8rYqo7AxF80mrh6M9yk4JouMjvY2+SxmItq098yd1GRlCbZERkjqOlXy+iHKa69G4ru
OKbnyBXkg7twnV+V7Ptf3OTyWm/W12fYP4bRJR/cXOQnywg4TPhsWrkV95bnYr8Iej4OW/zv0+9L
NNS8bslZ9Fb6VGx+wjnkHjZRIxfixYxUiyeAC5G7l/+VeVwWCakQHHuD1OsTnlb9M9AcXWbR5AKc
Zuz6H1Wi9EC0T9tBcC44wseHw84pvUMVrauAEaM4REFDED7fJeIhxSNGg6YqXbAK8OI+671u5m6V
D+BxTKg1ZleAxd1wqybZmbXhscEknUr9P0Y553qMLQZt/aXMbCXLLcKMxqVel8KbgtBgloZrC1l6
cIA9lqVFRVJyorKi1xtEnOd2iqYRhZT/RPBGTd66ApFOA6Q/7O14kbyaH4is5ZokHcjG1fh/352G
OM7vfr1Ayf8eSEI7cFas0VhhDFeFGMSj4Hty314NgBE7UC5kJRbPmPiemkoRRne7WiHaQ+qRF74U
r7LcqAiHtGzobk5Iecpy2NTRpqiHYyP5medpLBd+9JcolEqi5Qack/GfdD4Mz9bFRa6QtteGpQjB
1HaXhhBXJY4fJ0Rp3uhJgxlH8E8njNuyERfhPU0HY9tIyo8LBfXS8oR22Gw5DyvP9CiA088zmACD
N2Yf6l6hvlXYeUj8CXni4YTdWPF7scZ2S1LMwA4YsVnoniTngmC7/6AZlXO2x/ar5WHYIeIM0yTZ
zJwz46k382S7ylots+oJ06fdxfytcP0Ye9F5ZtYLVz3u0ZobBnQ67rSy2nHqx/rkhVurIQ2h62ux
bZI6v/TXcsJQqNDtx54iNpdKffwb0sDxNXI1CmyZ6r1JwGFEl1I3OzPzrncgaxz6A7s+MKG1v2ow
dq5vynMC6hOklguZo2A+yJ19ZK/AWpdEMThgN0jKX5y3qTyoInH2ex0C329gvMa1N9awc+7OFYSl
o9qF4c92WpYy6Eim1gFCf6grBn4MhbcTwpmtzezRXLoZS+B86w2qOjIhIt6ySBr3v1/5N9Jj2m4L
f0/yVfNp0jZfGU3mddjC64YOgiMySxwTQZnqvwYT0Q2O8K+h/BMc8pjdHIMqB7QQ6SqmnypC4XLM
/TwYuMe6p63pXjZXfDbeQIpzun/XXVrLvx/ec2u7dUEt39psF+H9DnMk1Iw/5QbN16ZTauB1B07O
wTfpl8tTy13O45gy8DMDajYw/KXCt26sPyQB1lH7ZMcuTGZ3QB0HTLsXoR0taVfHOiS61pV6DZfZ
xJGz8IGa4Ynw8Z60YvckguBo4Mm0DfkkB4St0tRrirVdVGwyqnE3ElMKLDLzYArr+bGOUvA1zcBS
VUR2mqPMAZouc+YXZlBRMVQg1tBm5/SCJhfCT2a9xBjYucFQrsbjRGwZqfsJjI/OLQdrtoYKpmWD
HQT842Tdd3fxKM3LqYx8IdWi2ArMefPhnmaHjKlaB5Sueccpbh6Vc4Iz4YfTTvBq/X1x/ZGEHiTz
XbXOs12/sxf2OOBr3niULHIrXcA/suGwsC8bHDxi8VD/W2FjM8+N4HyWecZFfu3nxF+4BIYlxOJC
IIyVAqIX8tV/l400E6AaFyNyJyVENUaarxjHxEtv25M1UeIW8n064vIi4VgYdS4VMErWOIk6aDJi
yMkdu2pTjtDt3eForBwwZbnNkAUds3UPmLwVZ96BmfrGKs4nVYhL+9njbsJvYOhe6IesQ2hZkeNe
wHcTiHD3XOjHbb5Z/6hGCYPzEIn7i6T9rMsMZik9kqmVyE+r+vjP+Qqcl3vNVB22w3LqiA8SmWSX
V0mI2HII850+XZV55fNQSpff9FVyK3Sr7RDk3kldLJpy8dmQtXQh7qPACTJZH87D/nx+dAyAGR/P
HKeP+DudgK+H6A9RtkGwYRIQVQJkrAoyWD/krIaE9ue6jIa9ADldeJVZhTqT5PmAOs04pdkNIzrL
sQmrtuMzxPaIivWKx2fpl8RM7y4+xQBpU6BJIZlaH3wFZgBgQRzKdy3lC/UTlBpTRZE/VjgBO0l3
zngMiou1D/UPlbY4qo9ayBYwk8YIHt7AHfCDq+/l9h0Dk3EkaS0hJmf9unAH+4Gz15sFTItZUQFP
u/N/GYFE5CmpGnJtm4iyk5dU0V9DxMf/gOk6WPajYu7da0xXeNe+3GAEyoaMLyhFr2khY1yz/oEX
Q9uJY/m3Jooa/wxePQ6PcUFDCq6tg99vzEgB41cvT2e6yXHfMBqFUnCkwHilDVBS4JWNF34LoQYb
Nx1Hzv7XfAc8Wko41/MGns4OZyxdc8Juz8k6+sjTJmIYnuuuUhf+aVDDhJZwHW95WtY8lYlAQoxX
jL+3E1NdIMJrw+53kQFFkgBC+au1mfiUSA5reXmebk6PIuTs1A8uoZnnxZDQIHI4Jcr63MlqgTSP
PQNVS/cUCexNESZtyJq6wb4U2lh/OZvKlRI+SV8wXocsu1Eyu2vs32zL6WPBSsjhxTRUvVJf1a8i
bMok9rTIYw+yhze0/CzueeI/mrKA+g9OTP4+NtB6KQNFcQA/YxB/2ATGL6+oKONSwwXowbUuDTyj
HIysArAXg0vBRiv0qXb4BpVd6e4Aoln4zmcQMmCwAZrP0h8dbG7sGs8UwZ5ioWmzso+VIotHlu+1
dlo3yumZjU6fVnG6anDli8EkS5MO/18ZH9qDsHWD1SgI0JKxLFx8USDPHGtO62JLbf4ODYgF5tmj
eFixF2iBCqvIfel7ByY06u5bq3KHCUEfqb4DQN9uHRJdy0cKQbUj8yKAbTggzkd+NQI4YsKAqR21
uoBfmfq+pswMPpFTzKVJ5MZ3V9YAeN2CfQrG/QsxvEJ5LwMrTFTilJdsBYeiU5+mydjyXNWEQZEb
SeD8ScnVMwBVCjWFqTQFXNy5lIKWi+r3cZ72GsKD+7fnnN2XHOUX0FPoG+oOQYGl/F5d55HRyCTK
QnW2tiL7xp1HLw9b9eHe6Mpv7FUhxF+cY7Cg7sdg90fPF6EAqM5SvxH+J+hTQfcVvO3tJmjmjXEt
toyIpBYH++a40CdmuDyTtT+5Bg4IssZ4yfmfPUdKfJWwaNQdplUAuTal60SRzeHkR1kMIuikpIIG
kkNeeaGV4NLEXoLgyycX1MqOlQO/VtV/cOB+Bbc27Lw41cy8PD1Q2owaWLlAKESjImATjKHCk4PI
4sHz0T09bj4rS0xZWreWr1SwiN7JG9l9phr8s47byeqY2qAaKvF3Hf8wy7i0yaibzEEutcSXd5BC
PHif2u+y1MQpijnwsSUq18n+m4Ybq/yO7JItWLGqqLhONqX9tfcWKkVPw9dWKPlCyJdM82GeDp3z
YpXWAQpJZcX8FWkdrfslKYHaYMu2pttis4tDmuwz9LffRxKBq4jSH3+dLGdSTD17niqvcCS/L+zk
rFjIevmcaV1Emzf/CC18qmGdefCj0RUhL6iK40mrVgqI4W6hJckBXYQ+mmIocOkM54ScoQyFoxBK
IhXT7LOOZ2tO6xcAt9soL4l5OqwGtVNWtlImqVmn15VjFId/wjmB+9HpSfs91ELRDQaLOaLOR2GH
GETdGYyS72rTeadLeqDwZi8jEdv6MtZ4aj6//lJK+9xgzWezHzXKsBDpSw+plDuBMRjdTyRiBSjQ
ADQllnifqvrjKkbnkSE5Y1ExjvTTzdEoHzWeyITdptlCseLjQjCwYWGlEH4nzxInzkiRFdudSCsY
cYvydRjFQwseJnNs0BVcq0M4jR7TWXuweQwLOQW8MuqBA/twhzQgVkqrBskQ3Ts1+Yf48YTS9Qir
2cRWin0OkfjvYuBRDf+JMPhulsBlF3JNuyZxhASgvhEcRM7K5b40YFzETOmzMPx+7qzoxgxcpa1P
P0YpHQvDDcuMvA5dOjymcimUvulaCDcHfx4xFpkpOg7L/UDjJQHa+NaZxl5jnFAlMg8lC/1UMiEN
EYirgKxvd2bVYPJrIL105sqiLHNS70Tjj1DWdleARmA2eH8S8WC9aX4hPlgo6Gs3PW8D6Pv9rbP2
vtwhQYCPlubCFq4O9aNw1dbaPCABLplQ5K5wnwqTwngNuBV4u6MVyShVQz723eKmk5QnbJHG9fT3
hpovdXTYgZ6dn8ArhiQZCS7xRBrQ4wohgdx6aJKo8f21uOysjTQoRZFBtsUxUFU0B+atYW0Y9bwv
UNgX3+H4xIY39NDDfYrVm4Z6idqXLHF3swOeW8ktz4E0T9uxxKfsmy/MG6SihVTwYdqDBxSc5qRX
oNL80zD6L9tvswWU071MTSN/0PFnP6qJJ8PKf2J3PhR8mxp92wx8x78gbTzcl8sUEUv9qFSizqt7
kJK25njyBISA9eJHe9M/PyKlXdsub5+Y/BsJ/ysFC4K8OoCJO29LF70BMLMh6fKIxS6E3hxnSqTP
NJmXoFo8ZzGgIoSB+Or6OMIyeiUD8HQkO5AOAkvNlG33msAlgcd/DQAOgE5b934ov8TzkWvtULoZ
+kQFbSLNihQWQymb+7jhq9B4cdw4K78KmfaGopp/KXgUqHT2ummN4LlPts1Civ4BY5yaa3ZmC0JC
zRtipt0xybwWodQUF4IaEA99yGefV0YfirRY2yVnjGIQ+w9LFJwj4klKau1xApsH5vpDNR+DX8qn
D8i3QsxAAIYbX+T8Ao7ybvpNFw8EbGLByEPN6/iPGCZpRkXaDU5PunLmQrhuk8+O1ygWlvRXmmNg
ybVZne5QrB+IrHoBuPXp8rbeCaC9N6ea4J0LzhoF+pzlsRLt1GDnq1EBH3wHWjyAgLuWJZsEtYOj
0R1jdVWtq2DJnyhvwFm2sCbZzdnyFQVrzHYc9duG627TNNJ8pEcaMAzVDQAK8lWAYNwg+uY0cYNo
emFdWEaCSpO9efk2tJHNkiFb9EHNWf5rlJBqHln2w0v61mkhnudKVcOG5YwdwnyKtjCEsRI96cqi
V1n5IHLV/Pn30Wd+zxCBIlBOIRAwQxsHTiIRWPkXfN/9r5MbkPyCR0PjOlRse0M4teiAOEKy/93T
6GQP4AxUvlanFGw1ow4a8jwDTeAsDNEecO0O9hGp+lsCHuenoLgcjeVH0S2uqf9+YpRl8VAcKf2n
MDXAMoHDzzMWF6iOHUh5AukKzhLqbuHQhIoUBwUmERdHDkUrHc+MmQH/2KHjKojMaGPPbRGGiBrw
Ry8PY8XOFzV8jT+lRVrcByz1bekE8YY9BjSx/OoJVejL4xYb/kZi9gZrYmhj6Eff5+fInvDuCH3h
mc4CMIGgM3nq7xUHiiJwGCuwcNZxgPnFkAIbLei/GKccGI4geRU7KqC8jf90FSt1TbKGhzGCDTT/
p/m7iMuYGr3HFnQM+evBvy+NsIJg7UWbeTsHPZRsNz2sWaNrmvg5KnjRncBS4Ph2PzTofK2sIVBj
gNfn8x94CSxyG4vQaU6Z2+uxXlrPjUdoPpl8ADw1bPo1dK5a15+kepkd7NEXrLnL20+hdUnPzrTU
+0X6Q/2DwPrtnwvvN14I5OsqpSAPOOcfzRKuwNQ4kxnLVPVgXSiJUGLdFB/yAwOBN3AhxQ6Y5v36
hNOf2FncG4VugKTgml9SqLa3D6PPW5HzX5vyYlsxZjZyV+vPkNovONK/eUg6HOxzaYqjTMVUN8+N
u6mCQug6P+XaigtjjF3bI4nDvRxbauTcxSZC641MhcOISJ4ACE7X24dWmP6UsJU+AQuj7d0HjzjB
WN2R8awfUWjuoawrmmkdfodMhUXFAOfQmgaN90UbdnwcJJvT9W5b+s4BoswjnLALDlANQG/PdFQR
/gKPCAVanFQUVvYAypYnzAJLAzIdcsmOcRW/qtb3yJHiZmmoGUxsdDjMuSOT2jn1SUu33AMeYssV
CPczkZuFXBC4lUDOPiXItfymYqgP6JOiC2GlJoVsxijLmee+H8jkS1qOJdLTIJqa+IZ2FQ0iVA7u
4ERMvg8KUwkr+OJP+7p9ws7XYi/e77QvQ1S3Cybfd5QhsqYTsXfrYzSKFdWz/X6Lwq73JNOzqjV1
W3K0Nj/7xoqKsNTmj74PoB7S9HxDw0ZqvuRl8y7FJt00FG4CwUMuW4dsHWcavaHq978bUFq9ulSE
dh0VYhUlt8wXb7XrH+iNq9ok/MVMAxIKrZPaD44X2gmJDmglpFKDkEOOU7tjl+vA1ITLAeBuJ0nr
5lyMnUX0Ot5s2jg6pdJqs4yUgaGwpl6KqCxzs8RlgSMwI4XYoXinPpI8RW4fWxbQepmv/6BaCwZv
oTBxCI+lO3R+o5T134Lh9EgZLvnx6NOQaOlu2JC4nlNAbuT8tbqPtDFrIX8kiXkoPVFfFglSFWwQ
Pa9wo7iFr5gG7lBHkBA5dBsCJRL72fQP7elLAO9hPb7tBGpwl5qE+ZkZQlPjIApBer9yEeYV3yEb
j1pJPnQ9kz86FPTTFrvnWGA8UraYtLvsUR2/Xbc1gOHKHzmD/fX2oVP5NRpTqla6f8clX29hN/OY
VXjPHIp7e9h5JDcT/JkwA/WEq9GWnvTWMHnj42VNuzTA2Y+Fu4NY0W0jOnIDuPd7aLY9mtYW/yeA
PHjdVqh/MRuGzmJvcsGQpL12gz9hdz03uoOYTT3U7zjRSlxxmAvXlQny19CFx+uIllENoaCsTCkH
aZmRCs/55z6QNXxXwvnx5uaAC7Yde4cPayQieG7aGFQuN5emRM4jmaw+LWFDZOigkLN/Kl0ImE9Q
VLneoNCIhpcE7044t1nGpKm+bzBWFMLsbnGVp+TPv4HnW+A7KuhsiLp4lYTBfpbGRCBiFQeza71T
artCx7zMPVbXkpCQjZKSO5uoJ3ejFQq2T9bcWpnZUCAE0LpKbiuXP0l6zknAwapR8mvoq1+2plB7
VxGLYWkaJUA3anhddc3lkCqy3lAyb+IbkxQ9UgPOJ4sg6QkyWeL6IDnKJ7JOWVMUiKtEIlekpjpG
Q2onpNIRgyFxDdxWATR9PQdHyu0Z6mszoVnbyeP2FOYlaAnL1+tlKCeKJ824zdzFViK4klplPYWh
5UuYLrTACyOvLnU1kBMY46QSNKU6NFKmn654n2dyZmObPkCdK7zXOOa7F6Oo+Bass0VXx+wC9Xpb
ArMMlBjnWRTdhw/G0jAybdTwMKO1n+YxJwcep2UwjnQp8FuUU8YijAmzd5BGPbfXDz6ncmjqdUlW
GGxMixiPrfmlSwhuDUZc8qDEbKVAYuSWE5EgvUndpLTCxFCRcPnFwTNYl0FXcuH2/kuSRh9Zd9i2
eUDfjyww/lennLSpOzCaK2qYQoeOxvfzkgCNX6BK6/hEREpMQwQQNrw4jDEIQS/OFGhDEy0XwzxP
Dl9+ienyID0xEwTJUvfEglzJSHPSANKhyWrI/kkc3qn3nXGxzeXdBbBtBJXUH+eRaOcfpbzR9dsC
7B0HhmM8p45nz7zdR1nMdzc3bMS4ckxWbJ4o+I15cGlGfzsmr38niXhJwcck3H5Z+m6cdj1YiG+P
wN6Nc1KqCOBbqBS48WRHJXzSUbD3RuYsX/AdHsquRvAJOhAbPpJP8nhbRd49bZ4OYPjYtTdiiU+S
5EoZUMA/6coIreVSJ89It7osr40DXb7bw13d1oF9C0Bu94HGYFpSENIY/4JLlOL+yqmEzAjteksX
KHmStKVLY3PQYKv9RqWvLv38xhH8xucWnPcjcXe2Z59F2S4dr6+jK7mbZw+d4v+QYOStGzfkB6Fe
PT6N4EPw/do1IOFYU8qP6N/ZAIJC2Fbhm+YhDTlgB3MZR3TOWh1y1MjaeIhk9G6OJV2euUe7ipL6
YvVH+twGq0z/VOZvcLSKLKKBSQjYY8FPqk/4TpODhAm3FhQ6UMKD/kyAdVp+TSMgEjw5UGXXCIIT
0dDitQ1oDMFH/aKGe0VDQov5+1lcaxyvB+dp3GsmhNFkmCB2rANrHNAqQ3WN4WOouAiepS9tBwtY
sNaRKHm+RQHe96D8jaC93fchNXd+Pun8sjojlsxjdsGOWCnd348FrcAPNYm7zH6jmKxIg+sx31wL
anpY7vhcS6gs0ITjo7xCev0r9ZNQZhinZQTBmXXYqI0Ie9HscKrBGeURhsuVIQxlXPN02dH6wEzM
MayPWcS9HNVLvC6a31RTjruEqgAZhfahLyNMPFPsn9pTA9Q33aZs/TrfJE6Yyy1UJPedw+i62lkj
F68P7n7+aEEcxeEV9i5oImFBEHv4K897saXXoCDiACuC4DUp6WmBIkKUurc26uG07ihJf1FclWcs
kgO8rsEXmCmDHmGRHSqZ8bmhGfnIDmpJPMoqKO9wcIrfby5+6X1viH7DVwWBp4yv08iJ74ly6Jdg
DBlpRgqGjxw+mAkrayatzcRdq/CHDWKV4uX5wnwfQKTA6c4OE75PUCuy805S5minSDZgTZ70TXRt
/I4uVRXJAP0X6IzGs55a6es/X7xYxZWueg03hClgcZKRsv9T+q0t88XJzQOc8SgNrQDc3kzgf7Y4
rYK7HHKyLGA3cXH5szX4Q5QWK1kGZ2ti3zNZy/g8v0lwvzjUjOCmPbEG2+cQXQXTfRxfrFqwBE9H
YNCfd7YXq2d1+T1tfdnuoI8Km2huUV1FnCxOQjQNe/Qc+eH2CE3ERdPJoghS1seQdWPqWxDf52SV
35pJC7qv1DElIdfqsjGifPjXtP3LOTJR1zyX/rzglFHkFOE11ri7ES14u6qqUn01onVrYMJPbMQQ
YJxjxINUU3nDLLAERShrOh3aESkjtpMG6hDk/R5y3LFUDQ0EvKqxeu2whP/nutJHvmdHRaD//5Ie
5iIpROclY0FvRwfdBmgLaZrgK6tGjNexMkFrvnf6UpZFkE39lpGXYyTqKNMQmAoncSJ4LGw94OBO
VF7IoT/7fAsqIjJhe9X8lN4YZLp1/NsHI13r5ot31RBXG/rnOTmYfjnxlPzu4FOBtQosZhjzIcB1
pjMT60SPrmnnzPIHaEhsRGflm+vlors+HT13RTXT7DeaA63Lt5n6Kk9iap0Xs3T0knD0wZZ8qtpA
nTA4JFEJhfyWZgXXWBBfS1bKwtBITwbkVSkITWVVGyzYKl4xc4HLYbUdc4nqoYQCTZKhRJIzljJ/
nj8lKpwmNyvrvH86+AF4R3f9QbjVSKajJrb9uXikskD7S0FNpiGtbcLrBztAttAcQge+atjVnwPi
sckRQPCQb+x1cG5MFFp+MkmrgFdbNw4H5dCww8eI7bk5r5D/oBtghbQiA+vQP60GKxqUh0QJaXih
EnMFED+KiDfnpBMZRtJM185wEo1hIoavfEYf0ZPQQmFn/Ui+Aed3z0aZeBZ3djdW7HWBeb2sZQwV
FmWy3OW5fDRKQe2RUt+WtuzDYC9oA0PrQcx8B8jN9t9L7izkZpy1VHnYduEIMheVD8I5MZw7b3m9
ohebS3TJaIU7/AsLc9A6hPvZnoxGMIbqsuGugJnnMUJ5/n+MADRjNSsHQNioghXPVYzbeLmvdImh
2Bxqig+6qT+K0U6HoDr8IrD3G4iU7ZlK/mSYckVTMrqabTtPKQ7inEpJQ3NpCZ23U3sctxGjDDea
avXjoGWwFrwbvmHpzHeL9ElFKPg8z5lUE1CIFSAZgijK/foU72ohMUmtEVqMclyCuaJfLXT0q/Pd
14Q/jeY11BQxK/7XP7oroNBQIsjU5g0V+mj+RtQJbnhPSXcmJHz1i/HslQvFttPGrxOgCk3TW2h9
xW0OxuOfKFxNHQQR1NwT5gKjMxqOQmryPDHdIZIw81dvABsSk5zy5jFoHNYL68gIGZpWu0yE1qZ4
7PclSby7o4jRxlRXv5ophWUZbfqVzXRZt+kA62UY+x8T1HNaplltnezZwgNh5vKd8CApoNxDkTV7
QGiRgdh0oL+O8Yk7B2qBjEt2CVoaOlXBEjb12zqBGochJpfX+4SPVbuZ2GcdEBnQR4sXfQYZ6fXx
hNGXxCWBhtPpX384tM5Vi2dhksd4Bnl36WB+gNjW/kPPUkQtUkbzioYSP3DSw5G7891UsVNFz5Sp
tg7ltUin5AuVg8XO34hpYVek0RxLNs7A/gPQyQ4903mF9HYmkBjt1E2iwvf8Q5M7ol2aTDr/22Wm
5BLbMBoyzYvKqEXe3e4RklTJYZYdDlIjp/aUMNOjxqaxQO7BKRsTedkzRm8UYQOi/U73fxfSJf+b
9VStiyPRPqk9UlnJcAzNIU+pMhpKQK1HvYKc2XrJqpcYjKHt4MbbJ9t2S+kVq6JhyQirnB7xPZyz
lwjIaBNLvbzMLYqARkeIgxyK2rlaApUiGjkpwPE8gy93rCo6C9PUKuRXle1TWPeWSVyyZI8cYU3j
rIZuA8qayqg6F5qPDbfQeSZB0P7MW1wMegdFXwlayL8v82DiSZ/eZboYkckv4fUZiprtfccJNOgf
moPJyTINASGwE4G/DYfrFAnlhfNuTag7NzZTrLNaRs2t4MwI74GGp9QkIuZbq+CMwQ0xkyRX49TI
DB7JFrMErRxNF65W8nbyUA6qvpIuwCZhfPyQGBMNyrMsAXcH9WKHcYmQFkv5JJcyDngRvNEuY5a5
wGAR0fOwhaRkjYZ8irRiLI2dbFag480paAWkthH1InsKsBuGg0ecUarMh74J47ESSmRpAomxYpqD
SiSHSS7qXcHnlciKVPhJQooJvApUcMcglOT6VuhAOiQ6bEk4nX2zcJizkVT2ZMT1PelqX15T1MxE
H7XG/PoEECnKc4G4IZPnV6m3I/7YZ5hbEAwrTJ8cdIfcnMPyNpRsHljMaXCNEYgqSMVepncFwYNc
H1HcClfij3wquYZmzRsiBvnubMeqSBHoCswjMrkG3h52A0orlV/CY3Gi1k3Ia0PWbMgB+JDNsMtJ
hOWQyat2nlnubxKtbkr5K5O3ZD5v+Y7AstPRueqIPRtwzbq3yJGFqKKdC0nvErTXCu8+mwMOPfe2
22v/8/Obju5114UvC2+H8FOMP1TN1x6F8RDVXnGbvyBNhroPK6dVlESXk0Vz1I+yy0HDMaF+4fRM
hK+FI/4pR1mwoCSIr0u4XGiw2tVaHm76EuwOSyCUaNpTNoomGt+ywKiikzXKGsG0IpxtR4xzn3d5
U1OKjDPrxCQNCLny9FL39QpZi/F5K8EpuCsbZBlzYjjKTze/tj4FNNWg6Et9aR2h98wo1v6Uk4h5
47I5fdTtUFl6UywwBa+VL1VhtqvFWtPa+bmL+oChj9Qo+H78ztPcOo1ylM856Qw9OUH+OxGX7CKp
E6r8mK0Gw/M+TxjYFxsgBpn1XdAo3XEi9vRZAEL1+5z7ASwkgA3+UZgPtApPSgCgSy38dzYtwAan
36z7xzJv23Svg654UO7Cx9MJxqK4m6RMErduw+DgaNxHbr8N7pKleXSFLlH99SqdAztKMh8OEpLx
7/fMuKgeVM1a5QPKo82yHemBlyBqTs00qu2e40YsQWlINH1vLoX8ticTACtZ977BVfhhVYheYL65
VWv0aXVm1a0jYgLu923kVKldNB6rM87gdecibjL1SIoIwNKWfAS0uYCrCw6eGt+O9L5whZdREg7K
4xN6YIDh35m7WYySUo8cNmDNwwlimAITQRNlBUPAGfCTsGS+cHXSJnDZtNpmOiZZvUiK5bPdsOKT
sLCHFjviTj776nISnTyB94czHho9pQIndfxL0Q994Tz7wCnM5cHkYea5ycnuBVuwdm0zMSlRVfM6
SvxTV50Oy2r88gfNzvyeYy2ZJJubGibfN44Bhmuy1lifu1KetNrPBw2Z26ff66VywgpBAMc8zOC6
6EWoR5piqngMz2SS/S5WqgfOO3kz12lncXXr56V75a6ULd5Y5ocUtPCObaNj3vJwV5VeDTWYWOSP
nx5ocWZRyqsNuYVP3GZVWGCPJV04XwzdD2JOBaahWGEm0NmVJaxA5YNtGsZIRUAZ5wB4rXVzgr2A
33uZPw0SMRITPxQF21wqoG/1XVJihG0tfKTTzjrtPYYEJDZgPUsV4wlEDbQPwSxxBb6TAclci18g
e/1vsHhlvTFuBfSs6bYY95H5Sb9ZAHFW6Dv8LW7A/CfrbdbDkK8W4PiV6DQwmuyuiodSeWm6ADac
908ZoDH/bOetsBnz2Rran+p2Hv4VRGnxJoaaoCA0sdawuMbenYLFr2bv/3VtqfFfBGoWfJuqM8re
AeYkYFMLB7o/OasuELHEAEfB+pZEVSkqayD+3cYJl0mpEmbVe5SAtn/+7sxQHQLXcYg5pNzZHCEP
JxcwN9FAQV4P0hEQfqjDwTMw4al1R1Fo4feQIHF061Pvlkk4j7pugFY0y2FkynUuQXa5T0Q40b9n
Cr//kmq9jP4oRtxKvgx5UqV6afjBZn5JS3t8n/gYR2IHO04cWCWU6ATyhxsbaRLRgposGji9uF9c
om8RD+3syHm1m1CLWwPUadoAIfOBfVpLwEOmxeuK2xPR84kO6KrhJHk3ljvHAQhjEqrKDaaMW2l5
9UrhmEHzCxB/ZYwNBjj8A2pHy/t0yf/J4qwj/kOLfEjl9I0ruWxY11WH+58ccL0SrEELZoHM8omW
zZTcJa+iC3jEVpyBbYnu1+Y0onZsFMGAqQ6HGu83+oNiq5NaltIXLvd/Agrd8VGjFHLjxada6Lzl
kr/2NM1Ha9BDS6o7qqzYC2G3Q0Td1EsCv7HHkV36JDY97KKlUt7jRM4+NzO4wzveCyloBIyUwyx1
+HhsC/i2Ky8dBDcrgJa76sy/T+Re65FFMiV/9O4wKtAEVlIUQC3b1yjtXHQtZU66XPAUf4nbkqRd
EJgCaZjhYVR4colFFS8nvsGsCDwAkZ5xf5puQwXjLmBQDZskr2wnHleUiSiMZ6/d3bOuY/jKEfwA
Gvx+f+gZEj37Cq3R9FhOW/OxwJ/P9+3W96LOIcivPYi8PXyQyoisTuj+9WKukcntNEHjFVlPxjQj
Uwjs1IJ3NgH2pSfovzlR7R0g73/Z85J5yYRfI2esxe/xyauj9d5iDiSt64gt75fij+hsDxVWvOmF
1dxLKDtLRqUvgpIIOKtx9juigoz4zsOszYbZnFOLicQaWRSOlDr2RuX9awdqFE9e0w+MJxeCMSyN
ZTYC5w3tPOeBClCV9e67GqZYPegmHoWxsLaLPaWFKS4otyBEmM2w+mDuBr/6PTh72sgW2SAdcAzF
URivpP0rgobf/YuzoDrUOjsC9DgjzNCQ70u43VWH8LkZsT6yKoeCgR6paXtUD/cFruap8+kW3AFe
YuRbr0WI0mOvgac8q0z1gKCzdxIm37Yvptgok+MYcRrv5OOA4KS/aLONAmEYCrcr3aqN4e0dw+DS
WQPwVKjD93jtXuO8JOOSSQq+bQqskFjwTYR25iQrJSkl3wKX8Tkzf9U2EFE/PXto1RbGzdj3BXhD
09OhMpAl4qyVrk6m5hzvNCADAyBo3DIfJwLCvn8HM3RJl1KLIhR3E/vXVs7rRs8BTIJrRTMG0J/M
iIhtCGQS6nCbSCA8vMcM34VYT5ZhtIezC+ynC+rnF/8rOKm9CLUvlR8JUP9d9ErbIbAs2Ddh7oIj
KyZg4pBP9PaeNOJBReHPacjYrX3IAPlU+CXV0MgZAmFM8V2lbGA8mi1ddS/SksEuv21eFPKFZUYN
WBCT4u1h8BYsvLpiuG1qLigt0iZsobO0VWzqGTmMHuw5rrH4tz8J/cdke+nmzzUPykjKK+lTswhn
GyHJYFfye+thBvp5JmQCEmlqQ9U56WhlAhTrxEA39/OtzoZ/JDdYrQDPD6HCVl7+b3zE8/iAaPbE
Ar123YpY+YKBifx5I04/mkg5NIZfyqcAA1QswzRvB1IqJ60kv8bT9J6W/U1PGxxhYhSoeByPHGml
Co4+l6zMOC/NKthlJU3js1JuJ90CxEI6FFyc9vUMAFIenS/jeUMfvOuE+lEKxaZWagRXRobCdUcI
XWjfU9NJMT3/8ULhHnW/QgFR6J1rgw1KcmcSzkcixM0MfeIUfM/Ln5o2qhndojxoLijOY4cPivaY
lQD2p8sZUkLEG55AfSngqwobD7NAr0INkTG3Kunqxjlujx/ThLgwm4TL86t1rHh2wKOfTvHzU9oV
AW+7FYKoke/20/Y3+xwkxw4yLpBJ5ZPqXMGG7XYVIAL0naWMJS59VLXFqIBxVCHujQVbBDl0PyCr
alAiT4CRjtMtE2nzJeW8fvX6FK6ax1V1XMRxbvHwPSJ0r5yg+cTSxxRAOsde4OtHlv87ULEdWN+T
lOTA1lVvzHF3wfBdvfJbpsacPJRssSGQMGtktBS2nq6TG0qmMUwbjsJnPTpfFSd4xQ8jK+tZn5ei
8zssRBADDCRej1lakA6rvpAG3eroyFF4jJ8NFgdHqIzI1CO4tstTHyWdsVMfrmbTLFn4zNZm4YdG
ehWpMQRsrv+cbxj2jDTZPrZUbDf4fiD91RS9+QWnrWdcpUzP+o32TxvngAn7dC0kqnOQQ2LnvrKe
/Fyf+qmKJA4Djw5KhFuBOr8lb9YytNTQkamSow3eIkl1yKNmknuEoUZCZ96rZ0OjCnlwRutWFkHW
POPJfVqTO2/beUZX+vgomTewULAhXJdjLhTbpxz8CXU10lKEIEHOvAJlsSCZqfk/Xq5RK/0Jrvjw
21G/ycwO031ywoWlJevuzq1ajU7bHQJ7h8OF8rbA7vBPF33j0ZTFb0leYud+VSo18S/OsjNIOhoo
t6HkrIrwInuIaRqi9q7AX+b+MpW2UahADGCXnG8LRvuJKJ1n5zb6Z/F7c+bKl7HpOfZ1k5EQFE29
xncXbpJtKIwuud0tFB3eFiC7MuoFZUOZkeQFFo7UAxmzzp1fVjFG538ankCPjvcMFmFboqc/u2hR
YoAC13AzLEFjk7cYne51w6i2NyNW7b0E/QRkHyw4+ZKrdWqM54RrodLJakjGaEzMMHDUslUB9xG7
rtPIy5Pi77qgRYoVOzN4c4WsXFZTJWGZjG1xUV1s1uUD9KxgWqoeJ104i7awTgNut2KgRS3ye6eg
RGRWGO4SbzFWXEk/ZMP7ohm9upS4kNGIJu2vpB05/NxmhSYs2eCuRTDm8qjphwILSB5q7LWnncqb
WApXmKOqjCbtcyEtZM/FvPeiijmf4C/Rir81j98XhzZxbRU5gMiTmwzoFA2qKW3DR5zPj3P9VCP4
bjkDTrayq7TEoQt8nRAX9Oc8Jkh3f31H3W8X+rXBBuXg0cXRRECI9NawXEo1MM9a5kLwIS+y91z0
XzCwsXy51RPIDkokmKo5T/TQe4N6oT08ARIXFCNNvGoLu3Q5//adKCxunmjHbgd9G7GKzNxC7aGx
KVFJDL6EiEW+32tHuecOkppEyDGfVxnYNxlbwrnCLOaX/bPVYtpG6GDjHDzhNQG08zndEFpamb+j
9p9s58yYzX8tHg676E/erpM1DE+ipwEQs1Bnkcuj4p3JJKlgYZ/q4rAQ/AvIqWGyD0On3RPRLynf
NN+WpvnBFEzBek9f4LbcBdzNPj8370uhy+sKPM3Fuunxx43wpYnzDnbL5MZFJGS0ntEYM/cMIsJb
Dz1yQzlEQatFTlTtpH85KwaRZlPQbMCMMwdP8P/bs0wsTMjMUpQDB41Ugm53SwSi0/KxOcO/nMUH
CScgAOHjiWQDkpyO4qnzZyy9+rixhnTp424t+IcyhvIHQMKrmHkje05E7mIzwaci4ak7BIDbcDsO
3voyoddb18IGXGWoqxFx81lmCKVKFJv1ebVE7Hg/NIOQ1C+ABqsmt3hw2n7buHckK+xAzbBzYuFq
Rbv1kvyHJYLFmo05zzpxhvHT+19ETu/NSuXI9fIWSttb+PVwcd2izOSziNT1sIc4zZdI4zscQRIX
GD716/BxU1rCRQBMtl11z2ZT/1owTMFYfSHU4FWIsS4thgSA1q82YFMiGWHzcVeM7g2J4+uwrjb4
63W+xzW4rGbiXks62gAeOY2vXLMi8iZmiJ8Tb3HG5wZMJ9cOI1HQ1ocvKNEz7FiqHLWNab4w5q9L
jVcwWJi5EMBvcpSUZ8mnSKQLttF2Nl7RgVpMaG04QTlIhD6lqsSOBufK5OrfBXInppGJZuapBHHU
jF6JrZV0WiwfPYrn94p7Jipg52awyxtb3wdpfB7UHQyzohlCnko9vQmrD6QsHqEdEwgC33MDRNod
wOthFt/f2uVU/cHShv3KnWtEpdM6MWvJS1XMgKItM+gWIXhNAsA4WkAke1oLZ57kaYQ9ipFGRLn7
TBcKKNIJES/c8SQyNoqBoR318RbBsxY+X/HvotMsgbz3T5eUoEbGn1U/6c3P1X8PNATLg6S+kbde
cPC/Q/WhachNGLzw3/TW8LZ9hIOuU5z3R4+3SFAVpmBJQxMR54fZPHyYHiM1Yenp2euKdcnGG39y
wOT668/Nkw4XSHdPE9AODsG8jC0I7yXe7Z4Ej2Mv4jBWgWGSEPNDiVJSE5f/B6xDPBpKu7UONBJW
Dp81hB2DUd3VbXNLa5h2WaguyRARCoEjcK3L20P5BpS0oVFmanqAMmJjV96JTLi0BNSTCpxX/NDl
SwEprBKfhN/D1JKRMeZHsvmly/hcI2uryDbv8auJdvAfkkMVYt0q+wnreSsRlszLtKyaTp1dwu60
L60+JHjPSaaudbwUd17W/8FOX2rTdaIEbiKpvlqcmEX8TSmgQh/3jcwsf9DSNMRr1YOTCStejFpN
D0SoT8gpQyUKvtRR5IUIydsPMWHD7tU/5hBXfM1kC1FI+6iHHaSIpgdEIgP2jjfARB5NGAsMdozm
bENZkRNqicDkb3r7bF1dhlUze2ECt6eLrjzSjuJOKV1F4NXaTBD4JYMjzgwUZEsBgPeTJgf/fME5
4RdxWNxg3x4UhWG7jStX0lDghKaJrNxM5ALBeNSaFvdiYHy+npGXQJqhDuC8izxi46Gm4wDm/nit
ntNnechckNV6nxriV0iD7KDYdxuu5pDRJD9yEoc85Hwp7m9WNODhgW3iV0XnAWcW3yvSZ02XLTeq
/tYLEGGl0l8PHa634O4D2yqjuxXJAR8u9wMQGgUgg8bN20J4n8tHxEL7nN59fZEBOVPLeM6Ewbhx
XrXNq5/Dp8+9YMypzb8UJWR4xQ2frJL5aqnkNlUDq7TegtXh9WLRAdl6rc9kQiFc+tlvPtpOLSDV
AR6jp/c2lpSE9Bx3xC+VBnROb1dEOqYUWX4cWe61PO05qFxWvf6YyTPf4cBO0/QBIUMiM17HDLDO
8yHszelX9FEGGUByQf4E1ssNPiYERXrWZx9zjAXxrTs76ktClElDIAhZdmMyB1qZKH5m23Ifn9jm
Awdz8savq4/hjj+nW4rVa3pLl0B/Dv6vHMilfYFwrX7E3FCdefugNfgrGbJ7owzdffdBj6UgyCdM
EZ35zDPo92mLvwDKXY5o+fhr9k/58/p/RDFAJUPhO0yGzqaZpY15b38DK3CdxPK9gDnJDrqmR/2k
ZF9yfMrx0ZoN7g29SstWWYtviK0OIV1wpUZ/Bh52+tU2tKXDZaviTuW2+CwQ/GNTaYCBBYYOui6+
8XLpUI0f352DG3krmqOv9eWGpAFDqKtXOahjQuwBNP3PoEYq06iIcdV3+F/Xh+Vs3GQemBTtm/gw
GQq5dqFiGslTStkoBmDhwIIFxZTea4CNgE6GhoQdnfYYAWvAd4vnGakXYUs/ZRzK8Logipj5CJIL
vbNYxF62zBOdHeMFa3sVdWqHVVay/DG8b5zku7iEZM17IZdFHCI7ZrAQXMgAoqMAnhMNiGiLw9R4
l1z5cHKA4U6BVagGeQNKfV84k5eNawDmikiC0+4yEhLGm68+AHFqK4lvZ9j/u2avGO8SCGku5yQe
BRP5Gp3q1orxR65OJi+/wci1lR8HNTFCyPiazpxejQaI5qWz+Z514e7UUhsscZ/iIWAkBsIh93OB
I0vQEDGtXgOEqI4MmY3/srG1DZl8age/DOn4lJjrMjsA/sWKgUndYm7o1aB63isNZW+BDSJZI1CW
Tib5dmH5RTPFlfFuON23kMQt3sgRzRW+uLpFH+DcNWA6lPbnnRLCHw4n2RvEiewerzKKaiPCsTOL
V/JHBRqq7ZOAi1laOqriPc5L9zyXntul9ySmoJvXpanVmN3K3JhyZ5QmcExEs/b+Y6O2dsaM2tuA
gs/333WXzl7bczHinDDOANU44JkPFc/7gPuFJC+bHlyCbouKPqjkyWI2BLqLqZ8SLtnQOsIi+H/t
awK6SXiBymOx3lJOTQqfnLQHz/wRJx/aZUrP2s6jb+T7O3normzz6RLB1z3IqgGEinYmtsarHQRE
9vqlLG52Vmp0Z0LcHX9uisLGCV0O0W257pORVlgEi3yNgxOpletd8EKrMTwb43HkanUS9mTpJaO/
uE/m2iGg3HwwYH8H2bZoeXnD0OUcocFCPg4EfCF71JzWZ01tVvRetHylB08ORN6MedJCKhibTdEL
FodL6l8HUGVseaZJ/W9HR9g6fcunkck64AlX+zrwbYWkR/Il4lt9Qz5Ofj1gbtMP11N3NpNCHf3E
E1MLjdqpXuvGSW8W6bGGmUEaWN+vPaNo9AjTl9Xf8U2xaKS2v8WixANogV1sZF8w2PFbKkMGahcz
dIR8fJr+uz2968IuAIGR+gZOQ7b7Uk+BJN+c1Fp695XcmJy6dQiW+Q/TycBPDhkgn0ukUeK+WzEu
8gYuV1RR1V4bglBuZOJjuSVC46mrvY9rUcCdkcMYmhiebs52Pu5xXKuL/i3XiUQnHUH29CMwfrGx
AgLlQcaUoBqA/5gd1jz5V/8n8ygnx0afSfce7KxepCE7sTkmB8JJaoFewYd37UFmk8LGVFxYwmWJ
8ojl/OsGLnalTnBNGaafxFYc5Df+ApHLpapMvQtZ2uxj2VCqFXVSiXOboeqpUBwXskwSZ14ebti2
uUaV1A2mSXtkP+gXxyO+wGndErJ3GDEh9bMIOgHcYqHbHp/7IlJpdw27+jVmeINzz3hydiChEJcp
xSjbLwL17G6a3FIXKBaMqO6pnv/BYi0PfTbGIcmYWCyEEwqShYBikemhiddYn0i0RZN2QQEtJBP4
qt4dOb4Tn2/mZtyImJDby/1zs8vL4eM9aVOWrGKfoCEB7GeHQYIlbT2CrljQG7zodolTfnBiqNIt
C39+xbKLdHqx/EgnAkIn25ahcE8oCWyleQrKia3otHX+uHLN3oZFFYM1NqsfXH6xLmLxIHhbjpCK
6s1gDVAPGY+yhCdcUv/HfDT5+GNpkfCHc8dYZqZKDU4Ota3uSxJpmH5Ofak/6QgjDbbraTAeQwb6
R8l/MWHskIaGBwT2tMFTV63i8qqXlpMXb9zNBeVgv8OfYeckdWhSbxqGTyVdfwuviowKawamVB/1
vrnB+j+c+w18yDIUu1+wDqNSZrPFAVkW/jfTk1JRcXwZwlt4UAHCHU2BlYuBm/RsMyOQpjnyjPzp
/966++WP2abNx9FkZAlkfHoAgOSg4XLgcihvdxTlrl1LXAouXLMUwdBtSNa7AvZJL+UrS9NJ/4SP
mmD8c2IstBxmzSLaNTxatZeXAjNjxqNa0gVFF3k5D0slVOX4l7r5y9IzH8NA6mV5Z7yM9iK/MTVs
bB3aGeKt53QgQyp1HEijOIljFf7iNYu38dje1kY4015Zus94uGbUaPMhh/EECORq0cFF+yyGTOmp
cDL///605evv0Z1ashDPOTCcs3gidrNNZ9Ki9NHKLKZL3YtKyZFQFwOGQB5oy9/1sEAGosIIwsC8
fW7IbEnoJh9c7lJjvGz89VTs5h8KD0Ec69zonsilGbgHingWcQqIpJ21LpOY13Bw8sysTs7Lrq7i
FxMQpNd8CDQJxzPGt9MhB1qzHTwPXQSgUjQgGx5wpMUzkxkzulEaV3eZ2T44BQMbx3C+X3UqLSai
fZfPRsYh6tbG1w1g+UFKkIKGCdovKo9Y6UG5AfthmeYGvO/LYZL3OBpLF/GAFy2j28vTARM0IpDc
AWnLDZCUsT0jmM4ZniaTJ/CHMkN/Uju29gVzmayZMDgld0p/zQLPUaCF5C/LjDudh4HPNm/LRlDO
it5FGzerngoCyMzTtQjJ0OdsbnWqnzQwzvsUnm0hF1XKnHPk4P+Mth+R9GlZBVdx3Nk7htda3pRS
hSZizDq9ar01DVkswIgQH1vKP33LyTRivZ07untJ5tpXqTv5XefJl1xGEOc6iRfMmyxtYIWNpmHe
xlmJ4oeiM7ESNoXH5zXlckdv7sR5z0rumCynB+E9MjLUfr6/4k01a4LFM83xGKkUZqRfWqTaWszL
bZ+dncXL4coEkc3SGm1qRv8BJ6u4tHNzp+tbC0MCGxuUZlWru8ojdlWD9HV5X108nwpIot6SVOC8
o6d9b6yeu0PFxp7YkSte/wW4O0ogrBjC/PDqwIFjQSJX04uQN795UsTV8r/Aja/1xri4oFr+01rs
+Sqs/6TXKwSyAyfN0nhtABW9OGzXZSmkkuyV4eLP0/V7WGg5CeBeZgvyTRdR0IbKYGEREB8/F3k5
MAZXqMMcK4ifpFybJZ/mbFmReic+jXjytU5YhHbGkT72j7bWMNoC1+MAcBhi+BPVT2ehOXJApV6x
2jpYnpsbBkblCYYzKn1gmD2kd+yxcF6KAhe+O48uw1Unx97Eo31Izkh2Xrphb/qva7r+6n7wphA+
gL4ocqXuBblM/kuLBnJbY4DWqINWUyAPgobebmOcBlJxtIA7+9OAhHUOfjuqYooJ3/7GloCJM3Bu
DXagO8lq2T2GfX6a9NdGiMkPbtyRvSgeQ7SSlL4Fo/RgV5jjoSaVYaGqsTgXWXyraPn7f4LGhy9H
xVmofOvhJ14tvwQb7DhKPU9+Cp5vTdPVP4xyyCuV2Xfof3JKPNa0QQ0ffFQ/kaK64EINHUrq9yyy
sdJalKlJgAO1AEhvQ0aR21cBh1OA5AQ6fvhCUU30RA3ifLMVDkpIAHVesuSr6caA6neCymttidrG
CxIxCga87U4W4MbGXKpFoUYyrBZ6+qz3jd/RrH5QwZk5Sbeg9drq876nZ0ss4GWWi9Um061/gEKe
q9KGVko8ilbjrqU7YX+XP2ybCjWHPuV6MQyy9LkMvW+Jao7l8Ej6/f32mVB3lhIU4fcApAW9BkVE
cZF7oNMf9od+Zu0f8V7YIwJqL3ZTqc02p+Uf1S0jTLAKpa+G+JDwv1HBTu1PDUAe51biksyjYUKD
4a2Rg3l3YQ9EeKlrY+N3sWHuHgpQ0SbE8KgByEgSQ4fb3YboTmgbm3oYBmvG3S1qQlLIq166ksoo
zl/xAnHUfEDgun8DqeBj5z1YnMxACemjGLDTOw5WimodBAkFgvytVkJbnVi2OtQ88rGCVgQGx6Sy
UdeXixdYAxgNZTxqBi3uNJpm9pfC8aaHP2apnhA7CYn5Cq3ypM3+R3BBizGOLoaxZq0pHXaDXlkV
W8p8nfMcUvFnMarUWJcMs1uLX4PcEmQNBPsPMBl6cRn09X+XikLauzvDLtshSgC6KuWj1k3yk/HN
zuLFTC/nDh9YdtjwvZeZEJqpO+twZSFVdy0Ca8T+OgGv4SErsXnhfLJ32OGtH71H7srE3mlZieoj
6ro9CmpSFF6NkOWm32Of6TRUwrKxGlDgQLsAM1sIAGs4dzOSq93LEsbFeYUlMKfqKzsPQUDxeptk
appwq5OeqziOzw7H9xRX0CiWMp3WA2x6QWpclr9PBhrv1OdMComnqExQTWO5oBVJGEM5t2kWW+MR
Wp36BggZ/q3YlBX0dxGj2mnsaWQWM2zVkNZ0F1bHGRWCfFLGH10btQPnX/VqO4WoaxS0zmX3EVbc
03l8FOZw2S0R2u5kwwDrKAStC3q4Bc3nU70x1hfPHnTGuIPm7gfslwqgNZ80UOSYicW9R2pPqyaz
odgVWdEcczhPe/2P95/8yzq1bYtrv1cvGejlyNuuERFJ6vbDLQA7Rv4bUnEtAVjuQT9q8J0yfo3c
QX2ehDqrMMbT6j/VFv/YddIpr/MD2AY5ZQMxxwfmZyWrlEjJr47kjACOpqG9a/sC3QC0X1BePR6S
FsD43e2Gij2z1eScWQLewCrPegGH6JOa24kusf/2YHi53A4yO1PnhPyOiW4XLCPAExwUUPf2vMGR
NA2mmMPgKn9Josdpy+Aky7USa/wb0Z3vgdSRI50BOY2pKvcPbAYy+xIArQmv2wgDzUSxgl8GhGXR
Zsivs48M48ZmfoNSUNRfmcWRLZIOuMqdbuXEGkhFKWPuKwQh8WXXyzx+Ts62eJt0TCawP8ZwdrQ6
+hdIl12H+Q3dQucI1mnObkYheHA1Qmie5oJ3Mm/siWGeSNPApvNe8pEZEPeg91MvD1SIU+IdapA7
49Kvyx0YyNwnr3uJgHjVrEaPdN0gyYs3kjiwYFGJMPg5v2mVXL9NUOlPQf5gYRzwd4AMCxzMgmIx
qFyedygZ9iEOMTMRe5UAfl2xdjxwWYuezppxzxJmWfxEHiZsgN2e6TlMvD0ANZ6ZbCwRRdfCcecr
YA4cEfOoL6RX1sCfZ9SS/kdRjb1Tkg6uUR4gmznvpTOJwCUjHtduOrNiEEGR2JEAiJG6I1u6tP/s
ZxZT4rpEDRnP63HEs2V+ws1BcFTrYLWUBLXI+mvUjq/glykHoSLvxiM6+hRBK2W60CL/gtjLxt/H
H02diU95RI9Wjj1ezMJ6/cXASE6bPGejomwXQSCf2W1DJqBNz/jJcWBrSoiU7NvIvE3YOXrE5Xll
bOrDcfW7RdJuhoiHUBUYx6i2zVf6HkuGXcx+rluy/TGmkFjivwezuG9fhlJ86rfsQd7Xi8BgE58R
0pDzgXrrt/TDc6gA6NfylLP1coYqB85FbjLLg4ozD5d2S7J0lqjWvW0QFyEfe9DTwSw/AqdlfTgB
AA1tm4Pyn9COjZv5+qc1mYfQjkuFpbns8TOKvSpAvAn+G6TI2bb6r9X5u6+02X5WjA0a/Su9ayZ2
Ze9vF/wBltObuxGWk7qzTFh/QxcBfIvShYcWEXP+ztDG6kOLwxzyxzWhURDGqx2f9gfKdXRVvTcZ
HqmLkXe9cWM/9UhgiOMdMuQh+u6LPdbp68Wx9c9VZMcqPrCqkmUnO9E9hG6HxX/VyGxRtMegm0eb
/wDYisQonGJ/OYFP0cIVFbySm4VeZWGPAvYFnsfaFCJ5RlF4u0eZnv6sHZalC1dk/eXp6xp/cSW1
WpqCXk+6ii/LjzxQGxTpEMlCOfG7NsH2LSvQF4rBEM+t1AvcPDRmgs5/IdsTVsCbCTgPeE05WqLA
R8MzRpoMZlS369ZAmPG5vOzVMNKTAZADFcMHjV658LZmqBs5KeF3n1nTP2YtSqHZ7lCMdptV2WXU
REXck2sbGSrnlpSDrBWu3PPpqJ+/M3kGPFT75GQpEEwRagYjGq9y1yf8yEFSaUqxJo3M5e5L+w3x
oYYXaw2k8NTkYYiX7Q6I1CXzlpC53GSDZHSiMGZOxlpCVdXtOmajGaGmNhBySoSg0us+xlAGW6HL
uO7934GqLS/HDIZo/yB5uhg4/12UkOmBfWKgKOFdrzE8nb2RCVADeFFVwpVKEr5WI/YQZi+pl8iy
8z4Kh89cRavHtKNvvAQReDfQvo9VUiEQYiPnqT33preAZiqDNbbxp+S9neYAA9JCd9FjYS6LrSl0
DI8m5B8NYrZC49YDgmtiIhJYKltLlRPiugwpr+YwpWWb9K9o0u3HidpT48IEbkV1v1xQk8fhw6eD
xgsff7PKV3SlVnphlLY3DS04jmsPTJvYBfIKU4aL5PiAWx4dAcgjRYwxKr0OSfFpQCbe9HbN3Kw8
tOw0sT7a5ymEhAtSwuHvDHUr47aIX9UY7Vh/bu5FQKXZgqY1III5kBOMxvOhhcih5sQMDwwEV5Eq
Oxv2WWvnRMLvLULMS1P7ysWv3DQHO3RW0M6r7LkHARQ5VN3Ek3AcCMNGXsSn1L60aINY7sXB6mQ0
hyUlnEJ6piCFIkYzNXzUhES1UsHwWNlk4dvRjpYMVfzu7v13QxSOAX2gHiMVRpinlPAO0eqOvIrd
0RSyyA5mwR559hjREvzV/mN3RN9UVFyfe2oH5wN0MZMNehfaCca/i7kzpnH9dtFqm+8nEBv6uyrV
7whRchRF3RObDFkG5l3ibXjolsOkNzx0fkb6QGYIiAn0M8csi9VpOAU0SNFOA2OcvT3UrX+LP45z
fjxxW+o5WwYSnUKyo+ByvCRM6Xg6HJXyb7Jlkl7uJe1EDRVG0iAmSN0tUxJsqdt284NuhNsdgij/
Jhaezar0Ljkrc/A8UWvMTN01MCd1Qg7Vl0j6id46V5F8cnNiMxbSlg900R3C2aQ2WvtK9hI4/p1t
PyRSQpM/cyMCgjN6NRuJLSPpT1Bt12Uiqut9ZVOTTv2AMsRANEkm9IeB8MCJ9n8nJVvvX64jHeIA
IQxn2RINCNeekwn2b2aXCs5c9sJHNoTJaiPMOZwCjHJcZc6VEPWq31UupFkZnPqKKbMZQLRNjn80
AfYEwLdeGzoB7Km7UcyJvLXqRu2WJAZ6SBVkiN2qv5lJ/CYp5rd1quMjpmkxnjazezs3w1PXzOGB
SOjML3C+QDaGKCvf6NlPE5jwS9hmwm1zi5Bs3N8WlmUg6ROZbqFE2gszaEPol70isSlIffspUS0T
6FKtdb+D7fB16nR3X8+C/+0nd2WhDWirSq/qmzSW22vy8jIyVUFdkQX9qy+aRDWyczexyDpyUvpO
f0K9Z7DTbk0vywP/fMsDMTm+CgxPz3yc6xhqgL0HrZyujS31i8buw+lgzxsgAkGKrA5VqcV6f3Bm
ZXEMU+smQXXG9eLVotfNd2JYr2gjsz3DRY2uY8rrVYEtPO7E7OibnVQ+k7LWfJX/kxuCvbvfDGur
3aAuDNMfT6E3uU8L9bZRtyRr8XfUvf9QhHq0w2fcK98ttGq6gkQbS9iXH08d2xgvsgDqzIPWe7Vb
NauGlcxAAFCAT+vUeNYkI3RPSL7S6m5Fzhpn1KcB5NLcP3PhynD0MwmjognXrHxfYmsI7RZbNNiU
I5HfkL/FvjI0oywlqXSAgaq6S2C9uPlJgNolbUNdt6d/yc/zhEFHIn9zTbJXSUWqOZue4AusE2sF
sLeR4sAjoxng4bymWEFrpUqb+QBgMW6VFMWEmErvYhVQnnClgtZNRYshk2H4MMqsMLO9EETE/Zs0
0MyOvmteOi5xePWKGE793Tk4zJ2KZ8cSVE+9j4F1mfri4vc43LF343zKiEGzxo2L1uaYI5bvIuv5
lU95IkJ2RiKtr6/rzqcCJgNxPhUQiGb7DbkQorIDojS7iaWbJ0byPWIu0eXkx/xY3vJSgIoe6EaM
W4Bo9eqh23zPslbu8zbNNU2s8UcOgTgOBSP7u8xKhSjSYNaDqLwnx3HTvYfN44c1r3FunK2u8jlc
a9XMk3SstEuh2tRfeC91Sm4As3B+UpY+23Nla+4wrOC1+biD2WJYgJrkhtoMPtwsN3yjay6RLZ2X
62t/oLTlYLTEKnwo82d723ZxryUbErCjX8v75h6vHRatZBJqXExxy2ojiBtcKpwydx+Iv8MWmEPN
pD9ivLncg3ktUyOYX2JPOKwsujUuf2c6VIK07xdc2v7wYyKHyrmvX4cuxIT7nzTyWpzQWY4rIkUP
2M8tlz34jdaiV9Q1rl73eOIsexMnN1aXprTN0xlxHDeH2Fz2LnI7QGn70Uyr1qGycZ5IMCjlz3Xj
eC2pcwic8GKmHsm9YYounQrXPALdPHPH2nJ91GfxlEqrkQalmyVYZ1O6x3Bal+udG/NvqOQfR4Tj
x89fUKzqkRJERrd6nzdiRCSlC3u/kiMJxiR4PJRZuEkE1uf+wtWDAcyrkZyxWO5EJ34SLjWzxteE
KCv8A2RW+T6Uy/Ih5Bhgz+Sp8UDDJ0g2x5qwTrlCwo5lFwx+68+vxREWFHKa92RhpJ/y9hDs0iRJ
QdYrnZ25JpukrSZo67C2pb3cM0UCZf5yUn6peO840FpLt5+2gA3OFs9PNRJle4oiAkY+b/XsKuya
KTGSiTiPFXjBot7rfjkiszwdmAJEzL0ntO3rL8EBSR3gHyEZSVaBVgZ0xWP/XUCCaBgbqLaDx3Zv
LVbuyfqT2nkbySfmHgke4Z4woTUALYpxNvXPPmgXy9EimaqGOdihrI+EwjwghOqBRjmJMFITkKYz
z++Q9P6E6Ic1LMGl7G8wd+1oK3220WkIx0y4V0hWXkLaaybVTk4ybGGLWwUFsLFV3gl+FBQXRhBp
XyBTNySCt5d4MnFbGG01YOnxNm/zEK+MMFFrfoq2IdBVggSWAfdBClYAKkizBoZNm0EgjcXJplTB
aHrvOoklQL4KsDj7o2RqHVc7LaVY3eOD7UP7CkFr2zFBoeYANaF7EiXosqi1ogDgGxSPVCnnBkYV
zsmi5VXmVWMZd1bg5rh7X33d1R2b12iAkxZM0PPpAjM/18J9bu26ZYm0A4tEGtr6jcdr531FGZQH
yMtCbWSEJ8XRUQEmH2dSza3l4fN/ks8rK/3XIepC6yVWWXnZ4cfzawqRYQuyM3CiM6vVX4tDPTcm
LwTDKTSOmTaUWbA0ybA6JaTFNWcZ46iph30xnuXujTziMM7BpU2eoPNSUPYXslwuFHLm4QWiEfmj
l9+YFxptRoiYUX3E2mZTeZYW4tK2eMKtYqg25M7WXYepTUIC0Ejv9bPTgmb9Tk4e/hzbba3e37oi
Wqqx+uE441ndulw6q6FVoMFmiuunXJAYuH0t30kszVODQq+pt9+1vFdD09uDelyQoTV3rRHT0Wtz
U2VoczaPGqM7aQpgGWhOTQdwOEGgQEmtKdZawu2BZzasuXdGJfQpjMy5Y9rxhXQ21ZlaEDHOHvWG
9RsazQPqi+Ta7HSt7gBFIuZO8ISnfMeQPlGBEcioEN+ypT2847jRG8dRFa8Ho5MuaW3jOFiyuEFr
I6xWGQ6tTYvSqdB79vzY2XhSIxhynd2NCl26gstk6SenX6gZdnx+73o/B8NIDHH9DE5+lr0DQB7u
gNJRot6vRSO76bxDmy0zYRV2g7Apz+qYat4whN8pHKvU9oZm6ZiMk0qt2m073o+khAM8IfJMY33i
YmO81NRbw/ct6WDwFb5TL45OJv+GY6xOc4zVK7nLNh2SBhKveKHDpMEf+9njVce0ya3NNcuhPTwa
3CWVvu1+agfh8yEEOBuyRqRd8uO/NswUiqtrKvv8zrn2OeAyoIU1Y2UIA6OtN4vIPF1r7Kt9snDw
4azJxepWP+7mH/66uq82FMus63jcEinLsXAqiD0tJScD7FOv1kqJBhd1SgD0fmZK3ES9TlfeYShw
7fo3GYS+Vk/4NOFUmaN9lwJDLROj0qDD/QfGeBaZdWgCYLApCUvwaotSCpD45t+7HVq7iFvmAW2C
gvNWNBW+1EPTBbYCTCJhzprgj5Vobkgtb9lhNUBsTe00G2637Vc/aDD6dkvSYz6gDStBwwdtI5hQ
pow4ytp9cj6Ge9Jsum2q5onbOHyllTnvhL7hm4GuaKhr3MlpHW2AdChJmMjl3Yf6uIRtHmHCa7oA
GLTklk4dXnDLiHF0OwP1cKELxW12U2Qhwod2HerNYAluXHvVjC+jLreK2fm3SHHDchTrY+pQMq9l
8IbChbRHI4FN5PYkhIHZDvQs0NGnDfMf/AENRxr0ffdR6biUC/q1rK/6jH+XguPLngu0J433s7mh
L6Aju28n2jEpl59trGIY7dgkLSDOG4l6mj/R0qB3aTuGDKdBDNkcBdwdGoKM+eN8MSCPikBP8fDX
P6la4S8GpRLYOqi3Pg/XAUKP0wkKjh5CUdB7HOQlhZdOU0uYfks34i13zFkFWVeLVUIGSMR5W5LF
QEUgka6uLOF1Rve1WLzEnLoDPEKJqAyAFVezejZ0fLwFiY62AAJr+3+EmD0I9GA9ZS6YvbBUyXap
RN6FohDMIRHK8bqJXtup5xiDSelo6q704j+rIIcl+82rXeIUOjYqUJFFDh9DoSfFXH0uP0runICw
xSPrhvrXYZpkranqesiEn9CM81WU/Ez1rIzj94HuZSFnoC0rr7682DJZpfb7iiM+nCaEwD5nLuOn
wrazaXrYZkssJNwPG6JPnNq41rcO+KAmgh3fCMsMkvHyQpaeN8wusv1blUDYNvoACYMPTpDHL+tr
mOFCkHkdAvNxxwDh20SIF+cjgvQiML73B0tSQtZ/pUHoVKWpI1gZ2SMtnD0OsxdOHlqGjKWwAnJu
H4R51NnzNz+k/pysJXnTu9t5Xbcq1vy1V9XyJCtt7TfEubmZBerTkrwP1AueQ8K+fmGJcpUGT9Ig
Ol+wmS+KvVbAnAF0DVJS0Hcny2LxQ0MsSNROBc5qtjkhBgFzF5iwvVSRP4nCq86aaR3W7UDgM0Jz
3O/2NicLQ+R6NsFdPqKBaidH6pAEOjmULICZN9fr9LV89Z6Aud5aMh1gcYY1Y5+xZjsMCQlXn134
aNe2Pw+75aiuHguWuzJaFAY2EkkbuoYoNFritRnidE0ZTfvrQeYbY/mfrwtJRbv6nDsL/DfqOBFD
JDd2eRldvM/HWTpQw+pv2Trzt+PuO06Qdp0Hf7RAZ4lLVym6qOvliCMgUDAuMQreUW11rOqyx/U8
nXy7equ7RwJ3qtEtw9hfqNd4pxdbzarT5rHIYqdIvR22kkn4I7M/yC4qNJXpewRRAd22uCuqBOAa
7zj0dgimzGHtqy0oq7rK3w29MQEx4ASWmdkmvtegbPkP+JyXzLJNOxBFY73rLMu+Pch0LS43DQ/v
kpwKXKipcj/fEohcPHQ3YAWIEBuY4GhfSDgta0hxTb1aRfe7TU8KmE0ZbX/JZJ44X0tkrt/L9S+0
eNRwy5Uv+TnrRgBmrT7gvDVNVt3GZfW5/rZp367Ij2SvEZNoN9IlJeYbqeODwZoEjjvT/fPs+gEB
RhMBo5sesFb4fiCjcBxR+dVDR/uvorU//DkewGooVs99jgsp9MVe/wwhpUGkkosqFMzJEjfuqnGP
plCroHIP2sQPLHNhcOUTqQo4dLxW9kQhe6WhwxKQ9lsZv0muWraD4ryLGf8d7eD7+KOLQaxp7Xcv
emAgqL5A4FAvK8ntf86qp+FxGxUhIZotWFCZmgmkm0I5TzWx7FBsKA8Nlw7mjVTIrsXaisS+f86A
I6Ua88lGdlDF9ofL7Y1gJ1TlAXo89vz9gLcBdtyL4KyvZO/qWHxmRscCd1ateHi6iSFe0ZVF5cNq
zWYIGHWdPZl01IMRrqDhAryHum+iZ1DFUA1KGnRvtoLMRysETuhTNifZRRxX56y4yNhR+/gno+9C
a7Ajvrsw8Mz9MuCi+MNg4Attz8bAn2RZq5ExPdb2c9TkHi5L7dWdbPDvG+kPMRezRTOZVpJDvbbP
AY6tommUOf5mGXRwznXsRDqfFyH119NacO/JeuZDxumT0JgHE+i6myYaRmLhaWS4qnpo1J57LcPJ
och75mt8SpY66+xkCezdRYLl/loPCkrV/duNXExUJ/rGn2YscdMZdWdfrc5PohcGcy58K8Nqqgbi
K6souTnQUY6WDflkWaeZVBDd59dGWo92aEFbSxwZnrTYvjVbe2ADgHyDEocBXLYv8DwcBH6yVFJG
8uFDMfVkrmGnmRkkPn5r7L7q9ZM+982Af8B175R3dqpqyX6KsSdqkGs4ZSTxWMQlG74xgUMfdYtT
LgLyb19c/RtCEH3mmYFvTQwtP5Cp6zeWbVHUUhRXSkMrzmWZzgcZextCOZ82CdPN0WV7LhjDGMuO
0uiyFwGHobabafcNqVFxKNAu3ILmyZTLPhqUzbVlCZq1rXiHQlawBw0hyeiriDziv57DGvVXM8Nw
ezZWjeRFCwwLPLiwrVkUlNJe+XFc6gwIh9mhP4zY41oCJ/mJfLKG5JSnHmGcCSUu4qao0zpo6I3z
lJUxsJCwwqZpjU5+0SwwGrfFTawJ3W4zNGCZPFj8a6omRYqQRwT2TxM5gz1x6s3nTD6GKNy3Vt5n
xMY6zr14iGDbkjsObk1f8fhKXSEwYWGDRRzPAsNJkMeFFHk6ySQsRO/dAxOXLKnEOaGQbbzPVQjV
DglNZQbgC8ySeuS7N7zK1ooSiDONj+ZMmL0cX+8HlaeuIoGNsO5jmbJDPpvezhdF4ZnSsAyIspn/
2V8BgLiC1W4USBaEKt7Jn9TNyne/6pF/4TYLIInJ7qgy13ciq82AT15o31rGF3UDC/HNBpHUQAs0
nzZ0KKllfEOhQXR/AKrj8q7zzzeFu1zE8FGEzpjNqNrwhTRLVa3PiPZny5rnR+dszZpfY094LVNi
NXcXMAC/JIn+Td1/A729snN00pJSig337ZDhIGxaEphM9UfOsDcZ2lnFwJfKHYK9muvCQyxMPDqZ
uHeM5u450oQxo2n4Qi2g0P/EwRuVebnOoOe6g0Cox8oJwGp401WMm1Ow2AG9+h9yj2wOeR3aesaw
0cieFzXXVD4d1UmkO1akrYClhe3du8Ca/Ux1L4rSL/rwyN+O7vdsxb1tnWX4bD2XFCXt6NJh0K1U
y60F8FIgCDfgSJTV7kk7u/JJiNjlyPbo0vJNjJHv9J9QH6lNk8pTqr5KzvcIrWkdm3mB3u7pqPYv
Ae0Ofw+S7DJ/1mVT0fn9iSsInrpfgmapguHvZ493lzNgPlVYsiSs1K9TrewWUgtb0kOwRy5uGKX9
7LkxQSYr2m0BKTuGGlCj7pwy3j31HmN76C7fk1/i/AWnTlHBNPVy+jt9Rrqw24t4qbYVyNxoAn5j
AJvx9ag1kMqN2+lJ9kWXIq2oPWBgGw2V5Srf87N8UHu5BFgJijH2798LeLiv9ZRmuwMCG6xfYlmh
KTb3TiVrpmQiSHCNrY4hYWuUbS5rYETOHTVrWkXvsM2dd9MCvqVprytuTf3PX9TUMYbCEZjfKZ10
izs1nkAJtx3DPkcfuNs6HX+F6+BeFkU6hgEE9ptvARqM24LaA247TQdBeTu1dO25jnV1xbOxUpAD
uN9ozbzacjTTaCRvOb6c1/w4HbSoeRXZf23pZBEN/i1ALZQKlJMBvqubHZtZp4F9oKkpHTxMw4TH
0vk+8HAlOjrVVboxpGodocgLGnDF8CQeS+8VQUNrf1HnetWFmWcPwW3L9+FhCKF4bzmNcg6gqjJM
GdU8zZQibb9WEMW9bo7yc+BtjOhdlDnLdTjJ6CX0fL0MS6+Dth+2C43yTOTD97OFh8dZv2zntsIP
YZj2AKJYk2hvyHM4hxOF+cAlyC7wZxpSuHKZUdGCyt3hOSiQL85N5TxQePOgoQt1bVuV9S9MDAOI
gZm4OxdswVSW1mQKGJogLdMTlVBBDbocf5W9bUfQIMNCghk+Z6uAXUU7VGW0euRyvsI48LZCZYb3
XZ3QL3eFOz90hfL3iT4Cbk/NueESlYv9V+36Og99LMXfEg6SFcWlvbokPL6YKm4fjbPOz2yTmaoW
vhiA53hV2wOJ3niMBGSGArMSVW7FSdZ6pJiVGTKsBFqJgJT7JK8GRjJQSI5hy6tNuFqlysYB+7ZN
YlEu7F6cYcncWdSrO90Ce6aHVLRiIiWblvjvr4f4Wv8lHhBqiUbXbMy20FyD6a2zfsFYChEp07LY
xzhaD89kt7FJl3lR89GwWhjRyAvEEcrMas1+MS8yursZsg6Tz3V1AuT9s1ksefsGNoKEqEnERYSm
i1RZTGhTsimfTdui4kGFP/YfXX5+oPb+5RVdG7Ia30FsBOA4GTY9HD0uuRBK8VI50+niHQFbl+tZ
Prq/dmXeT60p07o+ox51HvfCo7uqleKRXgkxlaqYq1F3KITydPDYyP/ngNijXl82PuyuzKCEbplq
BHAN8FQ5HRbP+oC0yEEn2XdKtH5OoeQWaDimD31YfALDc+R0huQ/chk+XtvaaXNgDjBv8OMACjKq
bib5klkqCVUTt5ZMAC7us0zVi+h6AdeHwkIinHhZYLKf0aN+BBC9GKfRc2BlUAHoX/HQejLQ3qt6
Ch3/kXGoY9lxT+hFv18NxIxCe7k45KrALW6A9N0OUtDQeusaMkP6VC41Pz5xIdQyVAzTPiyj9B9/
458bLFk9OJnD8EozAQQ9SchhRBRnep4LXy8Yq1jsi6OV4Wn9PmEmIgIj1xEdvBljJq4iegB2MmwP
R7sTUh9//B69K4VwPWuiJnMaBrA9bS2om7JZS1t7pHKITfxAqNBXbuRcqEmVfXKsNYSJjp5oXKbZ
KQRG1hoZxDW+P3TXovL2APYTzO1QyGoEvVEo1GhW5pXRuz5VhrjC5NchhCxwzTG/rQqHqk1WtWbI
oRGMwFxrfNzkZzSJCAe6tqf6T6QyVmz256kX7nhgqv3k9jkQmgXE/igsPpGydotbhEe+4fvRPVrb
vh988k8IR+tbYmEe0BFiduVo1eFNVh9GH6yc5XRzyq71QF7nKM47X/cx1zyAjaBLfrneVJa1qJRn
CDhB/l7ErJmgn9gvAcRBeHG5PdvgDE675jlcRL+RIgo8dTf+iXSsT8/BxbxspSeasFQJ3AJmtnXs
LarLiA9tuRMNg1LNH4SvXSdCtrGa4JZ9ey4YzDbjxdSRGEUqENE4A2Pjf7TYUpU/Euw35kn1K+Z8
AIE6jyhIGnsB0NSUsITZBgPF2GIwzw3mta7DIrVxC22QsoO4lBSTE8ME+1I70EE9H2qWMXOAK9jp
FsI5HRBNgLQyTBEaqmXWnq+tUGaIt2br2bmvB6oVbfaCXW/Va7RES0wiq3fy1FzP5S0f7aePNUiD
BApv9jNzfiAn/rmaG8nhw6LCnGC40s+8FbXz5GOli5oO9GW7xo3wM1ekkltpo/SiaZ8HP17NSqs/
4TlBCk80f9UYgaOypbgkG1T5JCb69c8sJedOWq0C62A+Thb+LRN846sE9kIUozUxtdrzDhqlqweX
d5FNsz2y3ElYiALf2JOETQxaq3LrqQt+O4GgRi9gGx6vFYTvvTXwepW3HWgBxgxI3anUXZRR8Yzc
wyhBCaWbUn3WXzVhFtfMT6mVb076R/hoj/xUCbvx2u8fZVkcnHRKPeSzS5qSm+6IC1/N5MU6rqmQ
Dej46U66jMjeHbLRMWqt1J5EBaGuk9mFTYUoIQOlwviZAbySRrb6koM4wsqHBlcl7ySeLUQqhYAu
D4Y8fI1UA+UHj305N1k8qLDqETqEuClBrcdbiZKWyz8jZIFrgixzBlH7tH/evkRkj/K+IW2QISth
M97ot19lFdXclQUXZPInkWjehf8L3mEr3x61uhvuWkDb6CgmgDez9/n65qCzqDvA7tQYs4vPE0+I
CNtUoXEV+x9s+4brbI3uSlZIPX3FaCmx/MhumeNRXZeRIAJk4ZHe1drg34931GajsWKW+1jjxRZ5
eiuZCCPfjER1vtpJIHFfvsPXJrlFjRtbvlepsc5xE1goMhthvUlwqX+OzpGSimSd312+ntkp8b2j
Gs0Zwm5LXVTfNPO1tl8bky9j7Dpt9OOZpZZwHL/rmQaozwSBw9dAmLXRjJUVfeIT4udPCUvhshrA
bNZldsmiyTkIhleuX62Il8PzYa7pPky8RKPTBmB51eZxg7h58AgdykvZJ8wXpVmydunHSYFFE7/D
NXAIjx5Jzv7KDFiPL4f3jggvAO6s+wt3G64AwBkLnqNchzxXoVqU+/vzv9mY+lW7WHMMyZOD5LDu
z4cTuhPgvZa+rpV443NEspDzAtBeinuzYDUp6rDkfo6FTApGME4tllEwFBlC96IlXO6Z59VdGdoN
3Ccg0TD+ihhFPwPPSYR2nzYaDVzJr5dPXhLZYySDUFjTcbqC9Qfhbt620wBnue51OoE+wXOTTYTI
M6AccpBh3hnHz6opN1dlz/HAmUwmOGcsFNdMSDiIv93kRwbH4ifoI1x+sRaMX/jP2NLIQ0KY8E4M
B0cPh9mJeRkXv59EkhEQVlNEPwkFr86zDj2XMGLtVOHRGD9UdsnKec5JyE+mf/EKdzy344MP58sf
DcTMx2MhjifTpwsuGoidrHTjXatgQ2+1tr2+FvleTA+dPChXBvCigQV3jgsFR4vRdO7ahzeTRamm
iMnoo28O/jaRpw0Ryi1wZSBZy9b9Lo8nWueDiwShn2qHELUp9m/PbjnCG07mTzYfM6aDx8guwIMu
Q8c0xEufe2J8uYNQVmWM+pvRj1DZix0wIlHPNLefZOcIzPYMFi96izLowvSpcmkYWMv1+chPfKki
jNwHQXA87cgpSDgUt3ZIOrC7UWBZ2N2XJTLaTky95Dy5EyespfSigLwDklvdRMsAO2F+cCmn1/Q8
EVFvDTj9wcr2WqnEwAESEqPyRA5gaQiV5ixymSZSTfrVhC9aegDUzSJUD1UQpmizbOUpgMnwxgBG
E1xiWJrryZ3wXQczR7iL3HaabCoWKAGB3aIsWthHaAXs2+0VEMEqBq7u7IyU85aiSyN7Um4rFxAP
9nfKEV8L32TVXaoIds/OgU+VKocigdW9x6jHJ+WWsrwBO9WfSyZQ17Ve+SxqnlUbNd1yThGD31gs
sjQ/vL8kZ01C1LgtGGX5sxqvMnU5brT7vd/IvvPHL972lREZdcNJvasIzlcdlEdJngonrC2xTi+4
r2E/H9uyNaND9cQVT48QbyWTjAqzIyh0qmQxDoUy3gM/pbUy9TsRIEMKvjU4piEljNEoE3Mlw2EX
i4cVZTL8vtbBKVmzIDjX5B9SAMxxXWw+ctki0q4nk36Xt4DqElugMRgwGgE7lFyCISs8oxIEZDZh
Sdn7Aq1b0/HW8DG+Gyg4mOpAnEY9isKnvT869+2pcTD/rCfck96dEytHVN3v4lw1LKWOHK+rREIo
RA+b3ntOipgYrS7hg9QJ7WFUl/Xy/sm+6OuIDH2Y0y422dwhc7ZPo21us7/3rcsoF+uDOviLDy0D
UHXGSUa0EEfmuo660n/YUKB8TY+A/qfMkaBO8CmQTNy/wnIf0SXin28q5oFcZgjQGAuBWKkzvpbX
R4Z8VTX32lBuM5O4uKSUJ0OpqbVLdRu+2rZfwcsaWxS+uwt7fQlKpeBUp/HRYiyIWiOmejDNCQTA
kgV8/epleeejo3is+sZVW68kikF5zg3qsJYOhy/eDPABcpaCV/CnxJkGAfU5jKeu/ltUoD9r5zs2
bzZ2TSLZuww+n0TR1fwucXBuGwD6TPZ6mYc+H/RUcgkYe93fup9bL9ZfZdreArJ3UVB5D0zZn7UG
mrUNBG7osCAnKk6wz65O3nTWnLrmbicpvlK41J+XHIkjG0y+BYMr9w2qh/50AhsRxCKJMv+3a5oa
7lgI/lW4aHcbozM4Seh1IkCGPgM2KBreklJgZV44fXGIsyDOhwl9SU2f2e/8nzhrmEYYnTl4RmYR
pxE6zv80mi5kZhl/Dabv6rtQRiwhPRU5y2cxyXc7My4qGJNpvGvJkb6cz/HFy9JTvw5S1vYutrhR
WsYPU2RJ+gVbRTV2UpJe5ah4DPg72PfwR5rknjSpUIQL3vnxD7kou1WpF83w6ZMEV7mZ9gdbl0hK
BAmqFDp611L27Afx7pq3qkupe0vgkEOIGmLcbwnSldKQqdGMjOpLE478T9D77cgWnwnqPG0sKelk
oBcAUsBxMhQEdgu0usSFGBXln/tMqKqlbL+X/Wu4DzANfNjazbbGo8YYvZySM3Fi3j+Plt6FK7e3
Mfzxw2UttYYXcnH0tHL+O9DtHnfr7AeipS/W8sSJ6PFJyvh9mUJKMnY1FkJi6YWKZgoTbcLtu//a
HkXyYe3GEQZZLO6/0flDnmYw81KsnOJcoAZadv0D86L28cvZnB8j/3f7xY1QRpPnndIzHFl9PusR
8ruSjfXuerzj30m7g3j2qRHPHZDRiu6dLGnJUQ548HE1Ahpf8B28hPPHDfUh60q5JaWW1VreYK+2
cS+ej1sO4DkBFRbN41+hUwoZPLKV/KZoAU4qDvRj1sJsfC2q2gFLW9IJyL2+meKe4PZKXy/qgA0A
Wge9hS2TcLHrbs86Bu3onbhd7GpQdNVFCGUpCzC+zBHGf2CUFkSxA26HEWTiRMasbRq3MsyIhnap
9ajFe3USY2KpCXXhf0LImMSICwiw03mEvwMaCDQTfzJPUI9ksxEGirSXDJvujpSbYPgPNcIRp/GS
9+AQn1DHveJT+hLjJx2xtNr7L7Jtt5YGzItU+eWFPflXHJovA1y6lTZrcpQjPLvA9hhajtlKmuJb
NVHlGT/rEg97s/33LI0QoBtPEJdHGVEbkpcnFNorPOFvBAZ3fNZoA7RZEs387jHscnHPMd5M1beR
bClHaJ4bjb/gNgonEFkVIJ91HEy2LaqMORKhivVvKrl5l3Ac1XzFYldpBGACaoSHTHDVRAJ8GxSA
vyMIyOyKLc+GZz6f9mwQJ7jyKy6NLIGql0H7nb4+VVLQfdOYn3rPVMy+27d/RtLu4v7IWqHvcfai
Y4zkt0SSNBCQ45Xqp2uhsO/CUQXZ0TgvFheYEXSV1qLrlOZNQ/VHn5CJ7OKoM0Audz3e7fI1T2w4
a1k/gEm3r3q4UudIvp16EXjiycWUihcj0AKvhR9Z3ZOwQfAtFNFBm5ZBGk+wB3/eAL4gn+ofpPX+
EdZ501AxnPzdamMunvk/Nl47nZ9PK4ALI377dX2lkfzJrsp1DqUrOCf91h8e9vUZPrvHDildE7sr
CTlBfJ4WxO2WLVoglUMO2kYjzzbzJWBfoar7oMDUt9VswULok2keBzC0aM5m3S7HLeAKdlqDzVqw
k/W9ioxJOeGCrw7ZhigGoRyDltVyLR3Gk5gD4PWVHKo0cfilZuqrGJ5kGTGZnS9hzAk+6eccWmtR
GMvhyF/uFeA5r4jNZ74uz5AryDxz1Uyt72GY89d6V3RfkpsMA+lKZCMSt1ebuJ23QjNFGgRQUgwo
O6GnQIvcO82RnHTiy985MwGAGx0qdh37J7TZl2K5+DxU5hsXnN5L5fNr0zuanrd3uHLUTREPamD/
la9pP5pYjtcEVfxTk2VTj7bcWVIxSNGYmWKgnNj00Bw44qfxK6+ym1SgRPd6IA+iDfwVSy8gEfZk
LwVPve8bwJMf4EWuvA0K7/+Ut8RHNRvE45cHXoNFfTfi5UuIbEup9t+RHX+lLumy0jJ17+U3m+et
leBQrA/ChZlNO6MRgWDAZ+QLyFZ4w5zL3iI+b5tjSTcbBpTVsuU8V3qZUwlb2oRRkUZjm4hGgnNL
EvPLc+euarNHs55bbZlG/oxABHr0qEiL7Shx5jBIlbwLd4yD/4uU+R1CJdceL9X4lrX2GzuUp9o+
vMjRNTsy8V2MtB6yVFvGA4D6xjmsU8P+udNPzUL/F/35isLjztOr0/D9Pr+Y5he0HkBS14TWJfst
5CegHMmpCkt7oDve3oOJixuctKTae996Sg91SnB+YHKG0zftU+3A8Px/i6FqSWIE2YpIflti3bB2
kTVGsNiXAmLwyEfrH4KNWNyIniuvq1szpN5TlY50vl/JWOg385qNXw2i0jB4usPxS4rc3OvQSpna
0F2+jncfOHBhmfKdsqNeTICDEHuEijTKkupfOrImB+8aB7muX+Xz0nbGWNVXDpo6DCTbjC0LSZiB
4KHBmMes5ozch317nCChF90BY9pTqThixNwZYkBfsoexMx5esi1HDynvMBZHJj/Ozx72B3BK04sR
ns7WIg5bYj4ZS8JUEv04GrtKL6FsSvDjadmpTBv+l+GDqJcCfEvvXzgxqaAQC/D5kfjEpcr7wQRe
a17pdVCq7lIvbfwLHwQ8uAZGDSjGzlkMhce1bvBsQoYNe1UHTJgEJfE26Gy4Xg5flBPVE/sP2Sq0
EHWlxrwvqAAZpoTnf45I7W/Xs3nR6ExI6wn4KkPDKmL5xwK8gORvri57uFxXRItXHjWDDRjViu5H
HOr4o1duB9VSWwuIG6N/wrxxXtNG3zE85BvAvMBiQxK/7kc5NTy+VMnUS2fD6jP1M88xlux+YF7v
zoZy3N2AXukdCh/MyfOOWDADCx7d1qbv+0vhR34wM9uOriNG9PON7WwM3qmRXIksZZyIRAy5xFeP
gmfPpvGPCLWQ9/RjhH6k3Rt5NdjIAJAQ+5PaoWu8aJU9Z5ZLKFx3tsl59ZDqjpmar4unRCl7yhyd
nel/iWOSszW2YP1WGLf/BT7IAyjWh1rBIK6H3kAQdDAFzSqSGcSJ/+JXhJ/+cBh9ePg/zEqgeMkR
RoaW0FMioyOicCgjWmoVHFNVW/hLV7Hs3qkdujTPdFZXSQJe4TGb4X1//KBmdv4RSyeb9IqtJJkK
2DsBQTm75oiW8k+9Qjfc4FWlTnFPQQzsD4iNjWIKx3jdNcidkPAy8MsWa6W+DSQlhIPW5ZO3VNTJ
/brAYexxI9kGIiRcAgctPFco1ErCqYSrGjGaCNvLGEasU0zio4yG7/xsy9D383Vc2oSY2QJatUas
lqtexO7+b5SAq1tC4agPjQUbMtIGnYMrz5lcsTSHxngYxZri7QVDRGGlml783JE9jr1IV2ItkdEe
Z7olYALmwiJnXuHh5sHVbAUJWDDTR7lLFx0Y2G6KgWPGGzMUXVKhil1UJ90QEjekTtp18XG2kf/a
AOa6TyrdcRFj94SzRSpvekXy6ZTPDzCm/TyxLOLnZpU6qvSC0supGyXtcNk0yksr5dC+ftm+/3fv
/QhEncempU2SLNqHreOQKvSESms4wgvjG6gFji/zI/nGcHrCWWLrmV9doO5Q9sVNpuVLNJzoL9qG
DYTAEHaPpagXKviy1NlllsuijMeJVEXiJMrG7rllSMyr6/HKditLgVaUCeeVdKCL+dfTK7ovlJY1
ss2IHC+gzdcl5JCAeUTNt4P3c6dwuI+hsWTcQlcrk+50dAGZVFm2fIz5h54it8pViKYf1p4w8uUo
OMjiQVo3GHybCWL55Adu9qTWV9J6bOHUjd1b411sB1aSMS+Dp6ofMZLrCV3HKn9f1uQk0kHVpEAf
UzypxmW1QUuaDqtRNtjMroLcRoY7JMG1ztr7KemBY0PvgnzkAqEl0uH4I87J9B7b2XGl5raeOBMa
sCtecegqj2+eG9IYOpZucNMvpXiUs6WkvKbIoFIWgumliLAuSD8OpHme4ieEnidzvzRjzDQsWIwG
rY2a8Z1kkpi0Ht4nU26SdP5+fOz8/j2NKjv+jqW/Yoxbz+ROdlYGpZlxTjuPFPg5RdAGK73bGKsL
CM/bm4mt91Qw00mNh/56PINzpp/f6WDZJUJyo91Pm4d+5mpsq1Unniks+h+TZ5zbJCuvyt57ElSj
61pLlYMZqA2EiZWK/IZs6wuzgRVXXwHPVJ/ETPD0WdujTwDYDIVOUsEhH1yCjCshzHGqHRoK/bU7
hFOF475uIZBfoCts1NXsNHA2vVUAFOWDx0LjxfrqT6zelRM8Ks+hTX5v1a9rndnT7tLwB7w0+8OX
pz52aTWb6Y62HGXFibsPRhmBo5RYe1dMZy+VbOkf5z/ypJX+okld9+oWyaTWNk2eHA3wr5qEh8vR
wQYRgb8FUQzkt9cgm+beu64g3PKhenfKxzrmvKDnGCkVMH9ASjOC4Ys30le4vfnASXVCpiECwNiZ
QVdvCbcRIqRFnwjHtdqBmH+EHk2vo0ZEapgspmOCbIIWMC93fRw6QnbbNVdbtf16VAvASJ6GSYDn
EsLqSATjbQ5YeYzvhKruVHyw4KL3gD6WmlpDK82Gh+DleMxNCQt5gJI9Tz4R8kZFbbkOaAb0OapH
qIHNZu7LfqUVU7SAEPh2X+TUW0L9zgmwUWLgXN8eW8m7tm2fkvSwPMzcr7W4UAAlMTxFTcT+jque
lmtRPVJC6WFxK5C4qD5yhezmCnX8tuXlmaVPAnfYKUO671t479ZU6ebCIcdoOlFBauo1tTdx2kr/
oW3qw+hZg3gjjwFqNKp9ilqq8oNeFO1Sy7HiDIcbM2bHKFSm1PMtjCfeLN9QLp8qMDGIpvNNG8yK
pQVqg38MLmDGqpk2uAnwHi+pCKWwMUBvvkw2gxpXi9ZLP8sLm/n73X2DdXvx3b0Y6s+hMH+SwWxl
MHQckcbkxVtSC4coKGcZCnefpFQKUp6jH5CZCn9NMoJgw6ielphXUf1e9sueLAcXo/16N+O0fmNT
Bovws0+/gCsqP9FqTWObd4Vjb9lA2y6YCmRxQ02o40G6pHifSUJfyaHg11Ogt8D7AcxrhBl2DA1z
D7YtUg+kKVoi875aDjFkjhzhzIUwxfZeG0+Q5vkkauxGJXM8EyyOb8tr2MA9nZcpo0KE1cCg4Uim
MwI2oW4lJaVPdxMwq6D4HaZfT106Rozf+cuugcYKbGOqJkanrzRRKnelTNnk+P7cYohzLjDlyULk
qCDWb0jf2z3AB92kRTmmIN6DylGcHNn6ANdoddFHhJFg4NAUmo8d1p85kROsfUoPSC19eQcjbRgo
a6QDq6YiBwVdJJggTvAZGpXcLQllPQkZxremdtApw9DE6QYzKIuDJv/ZqZsPwrlstUxheNRODI8C
faHil6m4Sm0OBFjJFFHxvKx8eeVCs5emCz5kZjhuBBfpS5x4S8YgyFP9GfRZN/nSwuRF0cx6jvN0
bWcEy7odaDd7csht2RnR7ZCnrB6J5ZaE5ArBJctRNlZdBAED8Vt091FCLajHMMTfJD3UwvMf28TD
9svNge/k1dgNSBg1uwT1Ol/kQX6JFbNVx1TeDyRmLXVxzD7FMWmioEcbrnAv4DLs13HYHn5Mw6Mx
Xtj+fR6UuwKrnKcx7MnLEZPfem4kXDkD0qK7CYFSye4i4sS3tRMNdcXiqjY4j47uwuCtvFjdplfJ
x4miAQU5X/2TaGci9JdymdLUVkp3bZk4ALVIeN/2GT+uaKS4q27y8dHHdIMc7IXCNFHytaQDXXiC
yT5wfpuAMoIBqf3esvrX/nMmitsltTmfULRT4qrHefnKOJXP7UxQX2xqYRaoXiVnrOgIbVhmUHrf
lBlvOVIT/oFkuxn02sErlM7wIPFe1uT135VSv5JXZuyS0rXjZLBr2sWxm2hJCS1MqVd5yM5Rc02P
H/nLl8CsNMadjuefFyJ1huYXhrcTek0CdeQy0SfQbgWXgOljA6E7KpiMgSXPVp2cOCvBvqFs1kG3
X3yGo89dwYHFUmCs5xw2H937nESRul92LOBSGn3/PNRHPmG9M4GtPioLMH1azlIMA/s7a75momOA
GICLQ1cJ5/l+3WIJ0bGfyRDuCFWvYrv/BVjjAM7Uip4KGJv/mCpGHSOB10AnZAMKA1cbAjE+HHli
0AUIDlBDd33SAJy3U+wh2J3OW/DLV/iQW4Z2JvJVgTWZ1CwPtWfs71167nUmkMCKEls9akBD878o
H2n5QEmEjEvQ4ihqNuXSll4US3esG6gMoy2DqtLUt+0Hg09CLGY2g34TDXythc/B6b2bNKEQhxhl
HuCYQv0J6hTwY0rbuO6MUdc+L04EgqA12yZI78pVr9Lze97D8ulG0qi6xD619gfCjL0HrlXnQ8L1
aGJXfxyB5LERi0LUHmXFCCZjigPBjqxnK5wi1d0TwTJIK//Cve2I18dOFvzC1Phmq5hvhFgau4Dc
KElyMt8d2dv3M4+xjLWhqNHY9tO38stlfjYmtSijx+mX2/6qQCmvPU112G3aQzBgh4xdQu3QWlLY
Y2nJ5R4TsXmfc92hZP/YuEP6Ees3OS8t567mqL7EkRyW/IqhSN3BFdHqXYcoyJjo3TD311lUfE8P
G0JzUzZJxrqVV3QQCtT9dhUXdLKVGg/re3m8y/mkmOJkCVaLACYQ1OgczS8nYmjBk0anxDff7qbo
2odEH1/qZBxwE1f7uxCWpP1RhHOu8tmab3Mp6swocXoYEtnzOCsL9mbs4sXWpiWV4dgXONOf0hjf
HjGGBurOJZD8TIiNJHWG8uZ4e1LVbciEF68uSl7pmpm8c13Z/ySowfXiqN2XMGGcyy4uSs6UzYg+
3K2+lsBcZbJJBylxMV4svaA979FGrv5UtJfIi3Nqw3irh8H3QqlwklhDsOaHY5bNfSVQgYn8oFSg
CbuMY8VFDKgDbF9SjbsK7LSI8Evi1Ln70xvCXPckLzocWnSuQ2xPOBOiV01oESi7L4cMPsbygDpw
EcsOb1MiHUbPlD7nfIkmExtqjQ6FAG1XymRpFsaKYoa9ZmyNRCCmF9mCazmKaqzh9++ZVtUz8wjr
8JGVygybnzTBzTinwIi8u13pXOuwx+PHqtry0Tc78bbzsv40wurK00Z0krFeRGf21k/Hi+h/Spdb
bue8JkbuZAKhNDgt8vwx1JgiZul3r7sgUlwqGvlKHwNR9aZoa1AZUIQiIuGi+NKXa71ejuda43fP
ocoq4Z4OyXdgIQPRc3SqT2U6WyhDIDUdFmlxLs+RAUgBDlEh52+8IGvXsjUYnI86tl8nImxKrPC4
/XA9pMFJCUKyL9N1SWN3wV0Ejj2bAuv2ovtgqou61kSw/zgSlAYdk+AefUMM1brvWxU1pKDfSc+g
6VWgtc80YikbN6KVCsDNl3z07lq84GfamgB+yFiysfQve+Oij2qaeOkkWivN3DSwwBeW+A/li8WS
jW1zvKBoxHAA7lGM/wCc7SJKPNC0h6RDisrNbX4FZYh3lA7FMLQ7bgdVw1y1HsdADDn5dBGeq+ZE
hsrAb+pJCieSpmX4aRTEirBwuh93jDUC+TLDmqkFYopcrAbL/SQL7KhMo+Gef9Q8Nu2Yr4BuTHR4
bUV0rmRym0ZnhMmvQwW0EQ79xV4J5SiczH4tMwBlWSwwwqWntPCMSQ8Up4TySAI0prMYAywP7BBe
kthDqj7xDnwTjfLXx0xmeae+i4r/WfdRbCUSev27V7Tih0tH/Icw69w6TjHw8ioaae8gksCM6l4M
shwB4QIqqeoUcVN4q5/QKp01yiLHoHPlY1WNoKVb3S87EN1ajWQL5gAFG3ZS/KO289xGGq6DY8v5
huZDRVa70PM4UhHtyTGo7WEMspCOs42U/YVb9XMnZg3KKBNPk0NRH8Uujdv7s0CA4lY35M2Vqp/X
uEVNaxb12kShw65QjjXJr7xb4DUeEZGMbgqsTRsltCMIZaLnZgirSTJpVDuT/o3QRXuO5ymCYZ9n
4qatmGo1mi2p2K+BcZPU+kqVwvZUCeX7S3mueBoHS8jkBw9qbaevk8wZdtRkm4fhcL9jPkA+AmfL
zQvKKvZX+a8uVB6ehjO4/JnzFZlQsZ7GgPuo/Wrm4eYJRk+ZA/2zeuCiOxOiomPtgFb12DIfxuCf
6TGDYEIlJOoYNYPHnDeToM4+ebemPahYsdoP4eNhrI+bIVmq6sFmvKphmxg4nG2s/v8pKZSMdwyG
NtY4QjgXoBYU30nYFb9sieaJjy1PGumyJj/YjbIF+2/AeljfKgyouO5lDfdP9LFrLR+g0/eZrbxX
vihIN88401mXJGPCYl6/4arah92Lodz8GPn8ckZeAGU52Yx+edS+WMBgGTnjNvN99vi9KvAK0NUv
NcO5zaFXPHN7PD+c0rCg/WY/piUtq2EIbUfJw0pX9yCXBIy30HF8860zwnjDkGs/8IzvMvFvE4tJ
07oRXq0Bot0ZQ/BhFcJLCSgmuKEtibVn8/mA0RTDhqarYaaidv9KFoc/PCPvqZu/92QeQJyAd+Lx
J3iVaBApbkOMZkISAemSBks9nDKiPTFpJKTX9K1qxHqoGuxJ1EJnKqdwd+TzAe9LfIlVJms6sdu7
BsHZUtmMsu0miVxDqWnQAuEuByQstjhxqIk5HWw6KTFvHg4nJAYZXhBBuQodRAXjkhPJxwZImNkV
9YeS6RdXX6BSi9YTXuFAd723Z6FSQh1V2crD4XxOcagX0WeWVjZ+3gXj4cLVp3NFLRTJWaI7GaF1
vvWUsp/3DWfrDrPofN2JfKLin6+5pRZWdmQ4v63vNRelgwpHrmJTuOXsXmNBnFPxhkKQX2XI/w3d
dh2B9wCccYuO2W4KSzxLRKa8kFGfeT9AfX5xhVQsK7RkwbUhzxTrXkzSzkniY4zK3+M0vFkR7ROM
k5ABR1spaubKO7YocuGiuNdaEJk49RxKVqkx5bdmKuuiXiDTLzh57FSEHcY3XWLzhbzrrcN0uZvQ
EDBe0mfv4ZNe6Iuz4IXCHboXrwuCbgUHVAjKsDb2jZbg1PUg2zJBhX1Wu/6HHpZg3Y3DyqXVgZHK
OCUQGNueCwVhdxQdKS2Y+J8h1zxlkbJobQA1a/UA9GMKnXl6mAtsSuKHDOTEKP0h+lEItv8T6ybH
Vk+tG/8k9cUsuoDz58E8qJoCAT1D8r0QPrHpwz13OHi0z1Lroa8vQeaNQvyVc0HuZS9QWxrZKvY0
k9NyCVHJbpVZPWhNcUGr309nKV3MCIOCY0SOZrJx1faAC2toyPr11RJEn5NDkaHDXoL7OfoIFZQA
iv5xknZZuk5Vzha2kl1O2+K6efRCtONYPphziGThOjFz2PnXSSr2cltovLPV+NFhw2SrYfuVFvqI
iTbI9i33RRoit0sulo6a6YHOhS/gSA6IY8YlMM+tP5tzrt/fCzoMmImD1+jDeJlT05yN7NQFCUxo
baAuqNcolCh7eVUj2tRSRzdfSom12Ss1bKmGLMZzW3JhOkOy7rl+jVOOZYU2VqH8GxQV9fpHx7YB
/kvVp1rCB3/jkVDJfA6HbRpe1wBkY6ozS45AzCn64FyEWP04fxFLkGNOwUutR0GCEaQfKdx13K2V
mEJGvXJMOQy6U//TsZ0ApCHe8bAVhQ2WE9oN0Lu8iCjHUjm0Ctls+IgUkbnDbGPhjYtGmRJuVxCz
jXRucIjPWUUQwfP20u1jMlnUKjaeQaOM8mgJfACLWECl6lfDEW3PRHbT/pZVcIZMhPQ2OxvgIwyy
vrMOwyluiLwSkTJF6lm1GPhfGNffSdvtcrp1/70lMN00Q00hYztECge2EsI+cjX8nlSaE3lf5wc+
vs06DNLAGPd8dhkaNM6YpVK1MOy3RmkjUMFEll7cwATJdOKweGMoBt1soVRZ2EjZUQzqEjv0MHPr
8yzcoCuSj29quGFYXqXJ13maeuu5iOlUJ3JfFMZMZVr2uPJrbX/ytapzkBdJA2BmEh8jeEucb5vn
wcgn8CXspSmop+04zCv5qsc6KOfT0QHrhO3QznVj3IqPFrgHjaVZvuHhYJwME1jZkZeSasfAju/1
ccnVk/DX0xs1L7uHoxPksWaLAQvhCG/Y2bxgfvR1Vcl81NYTFngkRqacXdUOOut6HazEzAin8GW3
4nRG2ktarPtoRFGlSpyPG9Mn+COyvhheLMTlggns2+ggCz/FT1+iOzWSZaKtr19Zp2JVn6c9WfnO
5CrBZl+2/DktM4pqZ5TRR5t/YLVvrHnFOVw0hIjULZU7bJuoEvwipvzPN5xL5k3d0r/tizmErlMx
jz8dNT7nCoEg4EZjn3nublFH+i4yXKzZwITL4+ElSeBATsgAdAzlANuFQUVmhbNUUKp/Tc/0X6J6
v8q/5DUlsZFmhbvPd/zOry25DwsXDyWvJoIcp9q+t58QEbpxgwovCYyC1K/LlAWJ1QIFhyeozuAs
O2Zkw+Q0GYL7+R9NKObfhGR2g2tmJi9jtHA+oF7KjvH4bvI98KdprDG3CeacP+sAmwXYfYAp5Q09
Zk3nhlWFEVg5qxEnp3bUOffZHmvSgR6VlCqugTRdkO1KqTZfIuEVlbSLOotrkMODYdZAH5JqAL7O
gTr1+H/Lr7SxRzURn+mIDPHXsK46xtnPtiKCLGI4UHj05JL/R3GzD6RTJ0vOkC/2loO51fIX7yFY
D2NUTTfZniwYiHfdUn6DT/yIDr4rL3dG2tiI7qi5EIyjXn2e2W6wpGrZa2MlnrLNECgGB5KcVMBc
oHlW6MRYdnZdMD0KFlekKxLUhx061I7XK2Wr/YNEmiAZgtGmUj98dbwnpbtbG+nY3jiSGdc5/vDC
sWTRDMrly7lepBbk2ETtCQZ62ljmp8uIOGjkb3kih+scfuo2SwoKDjnpMbURo9Ej7FMUqXXvOo5j
xVsptOR03gsumZTLDt6MEv4wOImIeMg+LwyZ1Ruao6j9bs8+NI6pJ8qAqWMO3DDlb5oDjw/u1M/N
cTZpEFb9233NXzjyOpKmmV0mYHfeSO3UcIiFE5QmNxqJ8AJpYajcy7IciUrpl7p7Bx7n3xgVetLI
c4QtcF5vco+k9QaEVADwtpsV8uHQoJNPvP4WAEx60bvsMtFAFUi8PNvWCxcejX4lVya6Iu3k6+54
wmfFaVhWa5fmlnty+Jn+HvDeZ+i/eS0s0FOqrj+9bxHJOHx9HykfcpjbHAKDxOLUHpq8kh+MjXf1
aeM2s7SKGIPsLQSwQ7QXztbWC5MJc27f1tUyoeH77nkaNA/zsIxdUjRpTHG2vmy48AjK4of/cjur
AZarf//mm+iFWCKv/TZ9cWOXoOpeTvt8WsuXapFXnAIqE8VOmj5xc90dUilx//g/0Xdaoi6ljriC
25YjeuK5Jri4mmKLDQ4cezEHulOPa/NXR+ppP7ed8Jis0SrhouktPzxoeoWbWlvbDx20S5tWS8D3
JVbnxY+95012Mf8xfqIlWEuU1fZJIs9dhz98zSocsdT4nyMoT5/iu0rte+ATkA3mT1Rj7xqJG+f7
x5gHDjTPw2o5FhHoBJrZnSuE6xqdi65Gi8/WpWWNIlSac6QBqim/h+/5DoOHSlAGGY0gBShJf/FT
5Ta/Gvzzm+bO9qgf4B0DDcTSX63hwURoJEYpnlg8twS9Ok/84Ni5fowjWe85pS0lhb3GrO8I5STH
U4Vn5u9FKW9R13JuoIOZqz58PRqRokaTTOPeQZ8cyBJ4kTNkLJGK1Fl4g9ladrtmaEE43TFhpa/Q
kLGqDFTFXgBOzyUERmDuJOJ5+rk8Y5AjXQYsdm/tgTEZFzkwNdDf5B7WMRa7HrEn6fWUQNVje3lr
aeT1eXUpC0TdvxXrD5foo5W76mAD3JF7NsoZqHfeL1opZ57Y7eGpl3AIQzIDcAxSkDP0pL1fAYmu
jrNr3+OWVtLSePrhXO8jT0pzUUzDbFO8uOulJZGyMneGLGXbB7gXpRBGxi+bC3NJEIWMkTphlLJD
f0wDWfL2BqOZwM5RmdC4wSCiCZJuhex4Pg2FjyHSLtUtCPBm01QJRUZ+F9Kp+E+uAwcGBOFTbqXR
k4Vq21kII4Urm1IqId+cKHe3fF6w+4CRNbwMkOd3gAYUUzGUBDxogFcG6ERN8Ou4QkawkI8rjE14
NNory5tYG+BdEWAH14cZh4o4KPuosTpAskTwc8n510b9eofI4SrNGeOTIqov2QDVwVRliUZQV4ly
jqkAGiKtF7HSN6bDQkb4HLdLcm7XJGI/XjvZriaWUgH5WqqGaK/1qmo19GbxMOoQzMz0ZpgwPV4X
SGK51b6oSlcqUdu/uughDWzlU6944ojBBHnmKROI/3gll1Yo8cMzNI8feyK4HSXjcdd1XQF42TNg
mLAY3m7tLqgAYClgCkLHQwCF42EXGdb/MItDjsZY4/zcaU7c+aq0rYAZr6ZDzcdZz1qyl050qR2s
owQMkLhzYNMfJxzkxoYvNtiUywaQtfVtndENeRiZSFxaE81G33h2OQ4hMOTGhBvqLWk82psDlcYz
mQxlxab6zSAL5lzNE/Lx6aNeKdUDbFs1pP+AC6rPYGZrK4E0usSxd7Js+Zn/6MB3+I2s/JINlMFV
5M+ggIJbFYLD/g4uS+PiT5qkNC56C5lVf9LQxKt13Y8Jdr2XfqsqhGgw3+NDMJbFOl/fiS4eAUsY
IjNjSQfbztwnkg88y3Xowu/63La8WW3gwD3FVClpYpdsXTTElVP9pnxyMhW0gpUkoQfPBiWsXSZj
knEIAtxrfJUlEDmbQS222iUpIT6Ku10F1JteDRo54l2kIpPobmfdCR67yXxTPhjyqbo4LWayvcFT
pN0VTf2DNLYC6CZ5RgfHCI8CTcK9skABeRvGxXfhdvfYEjBXEmuBu+f5bn2TrOxzHU50m4TBwg/k
ZzKzlWBORLFAn6WcrEyG7iEQNeq67r23EQ+vhuj7/TsmoPZrjryYL31TE8q38jI85eWueD6uAWNq
E/vrAnFLgbVWeStYDMc/s+C13QT70/vOQLOeMKRzuDe5ol+zHH8JKobXR2bji1d/34ehKA+RmqPw
8ixXa9cqVupqy3XE8PGFoadrsDxdDH1iwiWBkuNPX3dHwmR+ec3iYZM2yRmoVMfdZOFZWH38/pme
yykSwXEMuMXgUbGBa/hQZKdBIroOUqatUJYTa4AHDEqd2z3nTXuO8TPsMJI9tyzx9vmzWKwKmgvB
Dw1BRhqLKtvF59CuDdqZERXOzOcLQX4vqvDqCfPqQJndyuJ6q0NdLo7xXwxCKsYMq3ytztxZ5/ZX
oJTWZSzk1V+gqyGFmf+G6v6swHoOFkwqOTzD8KtNVeih+ZQoTarqfDsu33RaMayqmD5AwECLad7w
vcoVrbQEK8uSwBzYY2QIY5s9iXxFE0R1OtvIAm8V0omp5Ymy74+JYyQkDfFctXVIhLZ4i76eV8qd
ZnjYq9KzgK1TMGfOzDhLwRBpt5ZOac6PCMGWUvtxB9G81lsoRwTttTpLZ1ycnwW9DHZVztnYzPso
6hVCtv3BdAiuhBYB0pcmGSrXC4gTSBAhpmDAbDPlVCXvs58eMFhHbQzkLFXNnxFM+8AW1Ae+wNyg
6quvD3Zz9ks3YZVmhdr9nItld1SOqYmh4Dvchc3Sjbkpu0Vzx4I5hX6U9qL/GKVsHoNayszCVBRW
DbygmJhq1hb9TjzstcYF/97ZASrHT/w3Dublsqfl3yHf7LuEJBFqx4+AhuL/OWDZZAZwZ8j2KO22
GEFlW1HOgoFBz+klsVsfTovqcYx/u6sbBE7+nfF60PdyLewCdLH85xEQksUkmAqfw6eot4+SXgME
fQwzydtvSzydgaqw90ntFpqKn+0GZHEdTZfXs2zOXsUllU+it0wn7hJGWhDCwbbl02aSi0OfnAC+
J+rcXlvCNIq4Dpa/NHhskdiCZqUDciIiLxpYr3hu+SR3bWboRUMCULr8xF8fQ0z7eZiC2lyB4meT
kha27sN2j+GeDo11O7xkwXJR2DjoJLtyHmv+YG65uv5c8CaRf7eIYE6/bmit2R6gMCy7r81zOnGD
wBbWm6fqg3SQkqiG4ociV6DsPOcI5oulUGcVmdx6chnFA9VTlPAuzkiAYghC4uVsQN1J47bIv5+b
w0t6n1j3SIewpCoJmjeWflyweAE3qnlEZdi2CxwSX3xt7E4e0crBWgRLY+ejXhq1wK4EhDvDFmCu
ac4wVutI0sODeRaI8SQemnneUvqFWKPi0Zk2DiLokVT99xXWS0CX2UnZDIRqUXCNicEs0lOPXqYR
jtAFGCsUn+3YOCIzXAfidzYks9ZJ3LTdojwIEK5p63NyJahON6XcFjVj/FrXx6mZ04lfcKf5Vuic
5jKWboqqqtx4UhoXA3AzWOEYLziQl9sJmCr6uT4gOp/OqbIopF8Td8WAf2BHo1XDBA+IgTu/CWn8
/M74QzWiP6W8Pn9belVyRPlCWzKuSEFM2mKsYp2V8o9vyk+9PUzE8piEQ7x5oqNzW2vQRxLx+bFL
zmPV8Oga4DTYeD2Vx20lCGTI5No20i5ok5MkxaJVVeJAeQfA+/mFho8g+UVpK4LdPaRduuciL8kZ
qV4bLIoZ7QhONy2qSxxUIMus2nGhf6S9VRQLptzB77B2+KuRf4H6rbjWBZ9/7uIBXTbC9+efu8yh
bdC5bi39E++PmlFOhz3VqWFsVySQT4E6/e6NUcVWAJJGLhWn7ltGMODCG/BV1V52uOKL0BHzsNQl
h9xk7naJkjeu9k7Z3PCB6Htv5CxURdcu6WxIC3/QPimIDMjnzVAkTd4Cmb+77PeeoHfZTkhtaqbo
aJE6VuUEJOzSXnZ8qXSDPuhnnHPWDYoZwz3GZ2VgbD+qsxB6uPcQ+wIghu1QJS2pseVN++JcrTIM
/IT0cOu9tRhhXMrhP7TFA9sOHyKcmZNl8bnj49ygu2d0EOXhr+iAozksLWwFnu4sGv54hCWQM5ea
le+iSLiLf3ULcPchysttqF5Uc49M0GlL30XpNVlEkC9xVKtuvw6xBSGAOKxz8Av0r5W15t600giQ
aA3Ek7VEpW01oZAwVBqw8ZrixDKvKlAX8qEpMFQfKaXoCIyRkK/aOFbKf1feDZES7Aqy6foG92cp
ia9d1SoyL2t1M890X74urmQs/X80d4soKBmv+jfIP4WgxgSZdciaMWkbadKcdYOF/Kco+8PGdHXu
fxao8+PYB1SzyudXD6JPTf6DvaLGlKIvJCvA9wpC41MphuogwITQTuGSfStgiAOH78y+BdMtvASj
yvh3xK94pfMpZkN7ZEBr8tFA1KK/DcDBGJUQUrHKEr7uUbb4X+wjx2vdom/1p6y1u5gGhzKLhfIY
uQ+5iglcXkh9MjPDSkjr5sNhDKuQAL6p4KNkVoa4q1K7NdxWm49s4xNAlZnUcDw9QmDAGQTyL0IY
/v1gCJ6K2wVkLQtAzWzEUeGQma3XxvZZTBQ6pQf01SS0cBTDXrMNYJ3hRQbTUYfr5i5KswcTNpd4
wRMnhw8dOoOmKlNPE4EqGZTdfCop+R1oPpQu2mhOOt4LKHkRCFBrkYYCBbjzeF0Ce8yEH0ukIape
lVB59g88vnFo1S5jneVLm8xKoE09mkFMx3ucLx/12VGFhIA2QRFCR7E/KDnoEUw/Va/7L+05uJcE
MFEzeMH71kAr6TB/YDT3/G5AqyEFkVspMSk4Fql9UTVAnQNQMYq+ZUcF359XNCe8yjxCVH3/gDwz
FjfbOyF5kP14AzedQ/9GNJHSQE+tUBl99dEH2yQHanF1gCQabMxmdQEFxwEeiHIs5jhwUM7kHVSo
kOBTkPRom4wF3vdnursG82h9+2YKzsR4/67yalrKEcO0H/PjfV3Hf5vnTIOOFeLux/iOs+seH363
LfiQShGA+sPHW0jUWWvN1N0mxbt5RP8MC2PCHxKKDIo/Xh36C6MGadoYRMyF/NsjAYG/ndKmEHKv
5nYcE3284DbOsVZyyineQAz+zzwj5SRgnoB18tmhz9Ndjpyu/hLKdkCjXXzu4KrSAsNes2za8PPu
r3+amkX83JZusLCohl+NJxHX+cZJaIBKJ84EtP4UfE0zjzYbHuZnCo8rSjdeTeqE7PHe9uJKZhiu
IL690RwRiv37Fxc+9ItT+xB8vMRvwpKWWaycSQL6zlk+F5uWoJNOA/q1yckKGDvQgKXSUZsxBMhm
v6BKPVfiwuUMn8WBr7f3IihhEw72nWTJe9LPZ4xXeZtvmlg/4j4b8vYYL74PKRmo8ol6u1fpdj6J
KxyLdg8R4p/F5aORPPNjRARhU/PWXYmazg5yygJysdq0vjqn4HGyLle1A4A/AQKAM1ejMvfxH2Pq
rik6UN/CamGLuVmFsYDs6LXA2C2Qa52iSSEk0NyvjoEE8P8T3UXEnYqkx0kXzEl3Lwpt00ojmuVF
cOoDCyJ0hblVZyYb9E2/DJnjMaIp/GLnGWwvKk23fkG7TmjxdDeIhAqclJH5pKeGzdp04A0PmJNQ
TNBq27QmUR/jTXfxmB+ZJLfHOhYd6yo9fJSSahlXObaf4VaeMmriTw7GBAz3o1nIK+1yIaLJgsGo
mDlvzsxSos2YA7BpxdXQu7t6DFNhU8Ml9J+YS23AHwz8cexYZgO9d0vukHLJ7pEiBlUTyPsfukt8
UCJj0khYvGjWQ3kcU/6ek0/OJ69G49buu7+bvPs5sdGmM+XQy3TCdxajNKTFszqp8Z1rpIJFFEHZ
6xTdqXQssmVur0wnGvJKjV3ZaFz4P0c4GrPCmeckOCKGmdYVBfXaKsIune/vpHTqDocchU4v7ZxS
MalWs/0oiBKsauVuPGq2AaNNQ8vq+vHQBxrdEeEcczJodkMtmsv7MRflLCm6jbAFXKXQdxE4FM0P
11XIfeEhZV88H97itgZd+p8+z8UNjJ2uQJ4bg+Yc3aLi3bhKRBCPoKHFaUm3IsJmVX4NEjHxPAQm
+rcgl1DryNAlGU+I4FaCbvJ4TJ92Qf8xDN9l6jp3L/nn1PAHw6jYOvvrcgsNHhze1mQ6uCZFW6pj
yqP2+aSME84xIbWaYx+NnxMvEp3+BsJnxYfDMdfhQSOvuAQRidLz0rNoFBl4im8sHPP694J0Y9lm
g2WmWogoJ4mRrnXjT6gQPVpgj+2oDkLhHX7wE23zqYN90tN+k+9MezRK1PX84Ln+k+TPF/RjXEtY
DZAkyu19gFNINhX/jGuuWx3Dy1uZM1YyAtrFpYbTTa+OWEJJVDm7cKaO12pOOsi6BDNQaHnAZyZh
cJ9fTYS652miu/lbgGWgdlteUxaK1gMbalyYYD6pELKVS7BRaL5b5D2b/MOR4Hu18rzqsICQR4vu
DZTYTzd1YWwaQwMkmy8v/wfUxVDwGDSWTbgXTUrTuJ+01IjtTBPNxiY2tuLwuZX4ne72fWObURB5
4fbRgfVfSJmsQ9GmachnZorQfl3Gr+Gb2G7hDruurO+UDS4Q2PiFj4GxUzWj5gR3kpeKuG9OH3qk
lJo0DNmDrvVgIz/Irc4HK+r2FLIEHwk5CchoUqozkikid7m6NOcj6ktMRMw8jAXiyTAzTICpuAlg
7xwnIOxkfWXJ8InNfOwFDLF9Y6+TeXM3x9aCH7D/vkK0IK6E51E6we9x+oIBHBI/8SZ8WjsHFbtO
4SOsnKGCGrYQWuYwSh74kzrvLJtK1zAPWlQ3MUuGwmZa5Yxyp7GMlvy5y3SNXj+n9BPhL4TRyRo/
DFXFSfs8EVug/JPKKkgBgzDsqyn1zenjuJ2EOQY/1n1I6Ykf8Caocn1Z+BklT3CbUBGgnlDjZzaA
m1l8d+JlvCDP5v8WbE5ElZGjiGpcXYPJipPHiFMZaGHx4SslwP71LQQDYH3Ylyk95OxEFgXCYhFJ
HrAQuYdFc3mK62RYDp92p68NJon0M65iTofwl5XfZDpiYNsp+kciin0N5BVJUVjjBwkkaqd38nKy
0e6pjkH9F9ZCAF7ZdvPGOEUOGaFAhcrLyM3CbnjlSzlOVHDDd7BJ0RI0u/YGOtVhHTerqwo3I5f3
xsxi57dszvibj712oSiYAw++FhLQyJ+4ki5YFJKr7A/ugWsx2hd9MtaOyER5LD50dwXbBbioneK8
+caoPyjb4mhqfYUw3ZAEt2MFzHzkYs8z0SFOYqTt+jyZmXjQdNr5H70Jv/fsHZxL6h3YpF8pAHAp
fUvaT00h+LfDQeQbJ8UTCgcm8KtpDr5wBl5djhFPvScUgBAn+Ig44vLX4CIwyJ1i7Y+VjLnnQ+TU
t04OC3vNVkgAtNPqJdP/zsIm8bgBrlQe2sYlXuB1NIHLWX0/y9Uo1UQs4U6GJ0fZ6r17N7t6Ay8J
90vZUNwPqlhDnaHCBASY5Lm3AzclKjdAsGLW1P4Bl4H6dwovAGz7Tvr1c6Db6M8/HIY4eEJfRyWi
gf4Q/vOgMac5ftZttZA6WZV6jsc1oaeR0UPtAhYzIahmSzvUUWauk7oVyesQoVvf9NsLBMKaH9Z1
PvrzOPRC6wwB8fkIdGkPrBCo3uQJTZubeOt+z5kFx+Jnh4GkFAMqT2dVVIvySpjRqA6yYBexIbr5
gfk4nKVeW78CCZ6jPKjVXkWFRlz08AJrV9AbMBUSqA7rYl4K7u8iXmoh8iFxCE/VjdV8b3BntJ3O
7fJRhF1ZNB8LF+CmAT/YR1Ui6iKJkOVEe9BH/0jGfqA9S5ycuPWuqT/QEGO8e2nGBuXpGWYGChKb
HFOV5Ccy/pllljTgxuXySDM6DfEZNflmbNES00mm4GhEinET+z1iWpjqTQgE6+UoOq+Gbam1G9dB
cfl9WE18pwMiwkdwCZ9yKm7ysuQK9p9tNIRcuAGOxZuavy1vNnUkXBBYJJ0axmwBo/dbBNHbGpoQ
k7nWj1kqsFPBI+bG3hL1o+7i1r5Wum/bPriKMylEWYTb/mZOQXv6UFsoRNVz5YMn5GNe8g57zk3U
6jllPq8gLZIyKHZslEOI3+FG72qdKYWugltOUeRl2z8FI/nPlN7HmAblIv6+e3tHo0uVG9jwyPw0
cuxDekcvr6dz2N9nXo0ohXYCKYu2pW/J2EbAKUsjIxq368/eZ3UvypN5PJTT5AbOWAn9FLAKzz0T
j+iT5hEeLn4TDnr5Frv0q13r47E4u58/1KUw09RDZXHcyqPPJaddnFT1Y76K6Qteg5KQEu9tJXk2
CRvqoycxGk35Ujjm7hdl6HoMea2oTIwIvO+DmgeZPQztxtc22A/awh+UFMaJC2q+5s8mohDjFPNJ
HzwKcClMtM9cQrKT4/CXW0vXV9QdMhmIhPbQzO8l5xZ77Vw7Ym/9zrP5S547QQmxKIlGcKQ8yN6f
exrif7poUZZo/NHcrAQXztLS6GGrxydepn14RrFwY1Q2JytrKxnUSp1nFjuIU11Lzwxp4Z56E0Lw
+sZj41jpl5nH/5j70NhhwRBqxl0dLr0nT5toACmEreIhD0jGv0ys6NpgGHTMPjdqGuWPqPT4mJC4
rrfQuNvJfSxg1TikFr9QN0/2Hzi57utp0VjdYGKBl7dLcfSYFhHLZN6g+JQ1fhEL411dCABYhc1C
HxJnS6ePEOkXRKhaT+slTrKo/eSrv6gAj8vKro8XGhhAhf0ePMmDJZQNWxsVY/a9k1Y8633Myjs5
P6bFUEwIQn6muKQZZFSJKeHJIhURTad+2FajoF2Zch+KyXiFlPh2GbVLUzLLlgVWQP6i7JlxOJr1
6EvA8u5q7h2K6x1QqxbyEvlUGMlz+ut7OrBmV3/LJPGlHLE3pq1fJhKwKRm7cUyL25+LCCNpeb2+
pzUFXTxWlLXiXQy7gkwCnMMYCVRk8Lhfn6jR5ra8hMlbQljx+BFLTQtd7z5s7tU7lbZcmvYminUU
mGP3lEyyeid03W4h2tevl9Xb+72iPPv/gnazJfJLJWenNqTO7aV2Iyx6zIL0f0DmvOaG/oCqButv
6griYtErUt9+UUFEv6WoL/YTNJedQ/MbGPIP3b0O8nzanFz3J0GAzQsoasND1UrSJMbx4HDrVK/J
vG/Jip95PIs5VVBFf2f540PBvZQ0746eB5Prn3EFp591gab0mPJx8Z8EWdsTsmgZr6LuAALuzods
AuwbLBXuepLII3RUwZ7Ohh+yFAdIdxfTnVv5xhURIgmYAFAGtCehbdhsC5p87SC+te8lQaL/OYq4
k9ijYD1WVhSA6wolsM6VtNZp3aqKF8lP/8OaMgEUX93LFeeRmTDuOyQuHxVYPsbGDySfO1wMJZTE
/XOa4WXSgA3vf3ocuHoyDCGWPqLyKt2HKm3v557z6GQ0suMbY+0zjg14aDDI7XoFYmyVCqJrXjpL
hSR0xEsWyuoNej42yzb6wgrWl8Ixns5Ku7rEzqR5Ie+suaU22eRjzfO7FxRKMCxAhFN0t3r092Ht
jP5m/KAk3pI3HAfJUV6zHytK7keyzPytJy5l8Zm7YK1/oUaqIZcEglBiaTyFucayObi5NQeA3Hfw
ZKr1HXKrZuFe9/uXdDY/+NSlNld7re9xtRXOHm1I5GVgh1O9YqyzD/reN4wn+++IHO5sp7CDxDW5
0+CKnqWA8WmV3qhmDRznGWTl5VuMAc7O1C4/Y3TkFZxL66dGomhw0pEgz2u//vtXqXBcWu+b7A8n
+de6cZI3dfsW3xSxDWtdjcXVxWk9OMOtfqCh/FoZBw7tCpIAr+cPnoYJZp60nH3LNrxKO3XUrEnu
KlE2xSuFSnu/TDaeGP/8chnYS6l3rBeYSsKTUOcRLdB3mA3UcFsXkW9GRWYFvGTuLTOgU6TLRI8l
RNumyEzB3+SjhjDkZ6g0/4m6Lyt3GWtqXveLucZpeoVMXTPdiiV3IHQF3WWb2+JJ0xDajFEYdiZj
KLvm5P28xaar6wtL4lUPOo4w8aKtYc9HFPeeq8vMrPz77n9fPPx0fHENsqTKwMqyKx8FtrYh+4HP
ejGTjIn2im5kDAm9nhBw0P/zE60SA1JQKZHwTuc94jKqSMPqE6BITGiYYZMFt6Brik7Ixj1l0Ive
GV4GLsaHQAuNVe0NhY7IX9TD6MSAuz7wm34veueK1+6RFQm3sPNr3AmT85AN775RexZTGoUNfW1l
TfNrs7B/si7b5VNVvjbP/h1HKHfwkrF/hPGZ8wUShQWZhwtELfOCfzXJCWYlPysiW20sObBm8ZVe
+WS9j+8R++cRVt++v6GAHyzzW/b6h3hufPPZu/dWYSYxDlT9jdvxWB6Q10LS4t+tBMzQ3Sp229CL
Fg+bwIb+yj2CxNdwfRTwYqkv/3obTERBscSHEEW26lybUUx/jiZ40jPIZjMaS4027xXmfsXCzCBE
yQvyJiXpyOWcE1W4ddS1EbYR8QyVIZp3G38dcWVTkSCWCwUNjoB2eMV/PtOeRId5+xG3BwKPXG4E
LZcNNHUFruUaLezQCRgnJCa9XE5iut+6zoetw+c4qLqBLS66mWR/Wdz8CXhdX57/I5ZISXT3Rssy
f9aYfYDjfewdAIBArj5CtKl5C1Hd3lVJcRuHUkm5Zge2nWBs1wJrmPM0VQeAPS75AB4nvDMSOCK+
LqyDacR14E1hLP6HMstvjjJM2MS0xd0gAvUxXguRKD+vzW5bYHLOveRe/tRHgs2GwbKf1kbdrhyV
pAc/sIBEA85IKf/lhxuEL98Fo77yFGD214Ul9IEZ6RHv4M0Z83L5T3febMfDyeWEX/xwDoVsOyBU
mKK9PiO3On74WjPnZmyhwM3TNTcRhjTFXItr1hJ8erKgFZbMF4yzFTC2Mz2PTVozaVN90cUZgcZo
0CGP605gngoqoULNjDgf0qQoKDR1OoZYHv0pOMPQXqgZLn1RBzwPq9e4oDD0xvi/3j7LUlqSp0H7
4mu4h9OvhprnalhlyrKzjTzYLdtiydg9G2BuAryAD0YBwo9t7xWOP9o1BvOEnnv9qXa69vfNj521
ztc9aBl5iBuGwtGjUCaKI4Ybb+Wikc1xu4wag/UgqQvDwzlRPXtcUB0cwDBzcENxjjuk0/0tlroQ
ScexNMDBlSsX7gx37+k/K7HjaySzXM/o3zAECNGeXYTPPBxrHNNZJ1+bV8pm+yg+VlfT9Vpid/Hr
4HVv42nmOm9GkpBBwhp2r40jL/lIu0oA6zrAOruEFXUeS3P6wVoByYZQ6EAyDtPpdjki4mKmH4UO
MTGCWHqPJUjWeV1Z1X/5IASeDBgb4wKDzngjH5DBkXH5wd3ymdFdnMILNkgj3naBf2iNroXSUp9d
mE0ldCGAvC05WRY7Ces6MDLYqqY/D0b6WkSn5LUfhMEDnEccWx+BPQEh66ReJEFl5yFl/6+Pz1fb
YJwWUdS2HS1kLN9Kg8HFZA4gC4WtEKe877u9Rze6MIjvyjWZ7P+aHCpkLcdeDg8pNsYg6hSxlgqV
rx5GH4lM4Y8nAfkzefTUPQIQNMMFexQi47LyRyykuOIK9aFUUYaeekSpBX5nqZuTLPAKvludZPkp
ChGaW6GL/dZRPteXVn3sDBH3nQ+8k6nOvy+BBK8cBaHGOUyCU4C0l0I6yQqFMdGYC11q3NYhQAnl
/1sDtiCu0q/sBJvtHi9oIWKAdCQu4Xmoenj69l62FHOZd/eJrnPuR7BcQKWsRB5Ol1XmcKvDN9G2
kUY8KaeIA2BtUyCM1UCB/bpbD0CeXJjBWBbZ5j0Bu6Fj8zUeeCv2PtSGITtiRdSRW+NnNHSq35cW
5xNDb6a72hnUFDF2YBZg/2+G7ChIJr4xPuIdGN82q58QU69kkwj18D/Vy/PoPhevCSN7r2T/CoAp
bHqA629CyUplVhRTEkM0hJL3nkdm9LxsikeMf2PPmZWwvzh9OvEA7qNAgFpShFe6uF4iOrg6zPei
Y4/e5j+XHfRKeuoRab9Vf9Z0p53ZYDOxFl8VdIwWRSBUaDFLEn9RuywsvQWFwK1aHaLFsG5SF1jH
pnPumRQhiOE8li/i0YQMqqBnJxV0X/QZQrFduI+J4qEjzHuhkwCXvFTHF9DkkaC+3Ilev7vf/1Uf
hcAY3gIxAzTlcuCtLSpdxSCh/jLjeqQcl8HUaPWtNnPz6ywc3mep+VBrmKVqmfhxte6m8KOjiWOc
qPlffbEqN9GmTIuroqx7g5qCL692RMmkciKHFzZ4jVguLvyqV8nIozaKGSxEERLSJlJlN1j3BqMu
XN4vsO7Qsdi01xz/6JrA6HD4PbgPTtB6s0n5E/HzTo51VUnnvJIktS5vYOr0qbEqbYmHyUJMNdIn
Ll9IfNw6m0x5VU3AjX8uBXEQwhPjA7uhzUaKqfnMp8Knn5qYP1gFHVOmVJN8g0bBm2JfgN5TzYY8
6bUO6saqxZdhXAdUlGz2Hx9Tvo4MRvCl5smA4XeihNAHU6oCwJoKh6HN74Cu/oGnvvnywGHYP6IU
FbZ5JRf4+tA98KpKGuXwRKzZqkvzJm8bulpK2bXsOJzaypV71oslbhR//EKHG4nd7EiUXr4nP0eu
nbu23R3a2JwtcnL4909SNjdJzOc64olNIN5AOjLhnksd/SG2nseqREB3xfGyq07pUrePhp8qw1Eb
3VMSTITmtFV6WOSPGbICwwBzGcKziaPHHR6+lCOy9rUC2JN8LS/De4yYx+EB4dww4XBDYSzLuvKg
s0+5kNGqBzPKF/Yp9o9B8tC1KM+X2Hafn/z/TN3ugEwz59DdSRQyKegCbl9O9FdR17aNaBhxVK5E
vQLhGLj4m8oQ08XBS+raHAJlD69ePdd22LNHgsNPBvHHnuooH6t9n5u7n0EBjYGdlc67en4MutfL
7f2S1MySkyMregY+1klX4zj70owQU+icloovF+WGTx2aVAK6Bz+KlL3DbEvevDF7MCuI8D8FqM6N
1VyuOwc1v/rtfZVRK88Jhl/LbQQK/yddT2EonRbT3qHmn9tDMzuP8vfQSNuTv2Pzc/W+gntQSjtS
0GGfk4ldP2nQnBNYij1JtaZ7b1iQT+AUntksZQzOwCcBEnI0Dk5fnUledkTP6/6fotOrJ+Do+/Qf
MF167dmIn6qoE1zfUpMw9sEpcW7rY1lPMeYfEMEtvwko5CvsRu8VBkweCMnsBb0OQnNhWj5RdfCB
IofOBtVidt6vVZ40ef7fy9Icizk/W3R+f1sYrU38ThrsVtsxPE8u6I11dd4sCiz0FlBe7d2DWqgE
SWSEi6wXdBdxIK7+EaIjKfjWeoGeGPUQsPnBY/JGn3upjqeZmXjQNXhduk/ZLdfDBESQLlHqGxNd
b3kvNGz88ZDe/XySrqLgG586BetXEIut1aSCVbflO/ux+2dgJndRtzry+8ajmZCUQkD1Gm9hb6Dd
Uez7Ug3CP2GnvbOO105tNc31LsLoKqXteUy3F+3W6AClLJpamuJ57xidNwZ9bmfa5r2KVDyr4oNW
PKWZtZmYQE2m9Lp7/yaMstMY/1ylPvOmmVodwQ3HvOWuL1F/B/GFThSwgwdc5TbOHpVSi90IsNOQ
cekwqfluFfC/R6JQ/Om4aigt8AjVN5M0OHkQ6gn+aXNLI8+VleYJ+Pn3k0FKFyLAcdmq8sqLnyW2
i/ZrnL1IiY7vuEiw/m5ilKL0X1P9LjdXDnr2B0VijPLui0vteghKxYLKLY2NDTfvLjtjkZPkqZTU
/NbV0nisHn5Sc3MPRidbGqRMhUx9kf5sWD29gYgGoPAfzSeK4dUImDMgFGxLo98NAkQ8Z9q307SB
41w4/E4n8Bn0vw0cBMk53A5ctbI4oYzqFAeNKIe19LpGVTQx+/BF+ZfgSVlE3VxDrOmiIj7f7Hoz
MlLEnsEvPBfLU+FJeir87HJIcXT9n9KHgAHSebTwMlu7IYvF1i+1xgA61Y7TNojlVjdRwl+fHGVl
s8s4dNSwwnVLpQmwtlR5emeM7d8CQyqCNS5AiHIHxszQTIrwh+X3oBzGYAvyPUVSZVpY8q5Gvx/w
XRgHep08YZSGPUFC44rwERlwl0Om2XevtFfSnw2SXnl3cPlqnThJ1Pplp9MmZmQexXKR7rVrRSA4
K9l9NwEHqppu7FvUvQ4/jQQL4gt92UHHNQGAiZti1T6AVWigWF3YJsV7uKx3rlT6Og+3ld08FrhO
fCgVtbS8Y0DCH2RLSCFLYqqKKOUbDUCgk+3fn7kPIESqkKdUsY1YaXX6nDPd0o8suGtnMlC9snTX
J3I8NHQMS4GSf3NKXUN0xyJQd/YspvnZrw1aprqBSC4ftk4jZO2NqFO2EAtj6nosNDyUkDdsrEyK
CaoJ7ITC5IoID6m+OPLMwOS+XRCAIw0wESXZ7R3Z5IjH1P4lrdnixjsZ/QsVU8emBdiier3dAAzj
7kNMVg4im6vh+fJX4WgRBuPrixDcdIfMofpxNIjJV9pKVGBfOKgATF1qrYuKy031cRB567CQsRcg
Ew6W/TqbuCMxOTzWaj4A4MdnzrIPGe124Hq48wcNi22Mlpzzjd7wIMpI+IGlVFMQKD5opz7idSMe
nthl30dSyV/w9nBC6CEgh2jR1X7d9tHzv+OVcYvu2BHhqykoWU5uP+fK8oyorvFFPRDkmCboaY7x
ShLIkjCEYk7x9HcO3ua/xg8yvovW0ei/CtM1hu1/8jA1ofuffuU4wkPgxMizcJ3rxqo0fCUjlxym
qU2GzzzU32+kn0YY7Y6UnVJwcu4TdLGb9hQ5SggilpO8Hr40QA+/DWQhDlPfx4yMzuRxS8UsSIu1
o8HzCnMOI36z1Wpyg4lrpCfJSDp34Y6HXMB1kq02nWcZayZtDXY72QOncbXZzLkBKOqtWGNg+/OM
XENcQ/8ump9IMTl0uDNcNzhDaK6PglSPaTwVviXJUvP0j8QlyTG/UgW9G15bfe8SNR/OZE7/Gk4r
PRnuv+TBunpUg3ftpQEaFSHd8DDe2JPv3K5Xz9mvGiSe909fSwOrmpSigfJHLMK6vBLtJ+L4Wjnm
hZ/vY2RfEUXzs8/JO7DPPQEobr3ZaVwuffK5Un8pvh8lsuOMEikOPRcwD1jHvwcQzGfDMIcMhoVQ
qfpPqyy2PBBW8hdz3CnfQ3fq6W07iQH5mVxEXT1ilAwJqOUqQq+zhw7eDWBtji+xZu+cX3iicTYD
Wfo7z6VEl6x42LJt4wRtODz6423SzOkl6kmlcVL2fJNPCZP+ZPajSt5BZdCFQ0+gEkWbhvUHDvOW
FlHs0oIVbjnk1uZ2mdm2/8bZzfTjKB2FJG3J5XUAHwClgV6xStTLGvyde9z0DSelxGExcs1MVKTU
YrFJzTltw+0pbXynQsTaLje1WAgge+M3amAp1ZaqUvRfz9RgklBIGG15iuQhbc+o5qqQwvwb7quw
MBtZkjRKFMrPLR8cH/mveQ4f2biT1QeXPLbowNy9Ta7qRRY1eIZm/x2Z3JjvHhTeq21ji5aYzg8O
anzOhprETCt6aq/u1WZi/5sZRLlxMn+BUYUnjzMz4wHhKbaHF2syvtosOiKay17gSqptrx89YOPd
gmMNfb9mTQOTs6weiRhrZ3VQfdCo//k+4YNx9rvyQKbXNpT1HaTYXJtwdQw18SRLjPOkYBDv+l6U
2WCHV+PqLXhQeWXJjekHyhU7tOehStHXZaN1ilUMkTlnTfZm6gw1uPZSBoH8girSvFa5G7pknpPO
kWg4YbDXXZiM8uhFs4eX9bBjLHZotu/jfIv7+EJkoQnbuc5RwX1SwwPMxwr/xqEYeZdBOaidTASx
/ygqSKfFbYXYusdF5d8/lkJ7V/MoOCkIFn6E2WpA2BWPFP2j1gqXu3y6rZ2fQsU4Dxg+1L6CPzJ5
5QsvQ1xpzRs+EPRYFMXy+Kbp97WaIL1BHmIWCIFndk3Z6f1pj6fVuAAJKKqMtrjdC+CURQ3hPWxX
31IW/dsqaT/DMgK8WWaAm3994awtMpfzsLLlEt5Ww2bq5pLTwGMCcKFYYtBc41vhVxlKcwckGAsd
ltnabKx23axba9rYlOsYnRnCXPGl11BbGSVSp7EEllEn3KDTWk8sybqG5j3enAM7VtCBtJPt3+L1
8T9ot2zWjQY7eeIfUlGtR2ZbtNxCqUUOaajil5ics7vmVgH+sRMz6Yb3Ldm44vJxJ/pFCnzRMPlb
usyLsHQ7G4zeU5Oqga8pNQ+FjuFOL3004uNlq4UPNClm00gFo7KdwFIl8H8TGBF/i/QChX9lcIqb
rBDwDJpDZ5keteRVM6rP3TGO0FQNF92GfgWeQUfLaSweqleqyYs1Ra2zfmK/2JLwccq4KRNzA/6l
28jZO1XnJ0dzS1t0kP+4PRrRj9fCYoukxWRi22+JUNiqEPRW/FDdVUUPBJ57nDPU5H+epteb2Jmj
+YqAO/noNQA3IdN8T4vsT5w7t3TLntRoBk+d7F0gQrmi44L9f7qimn5UskfGFvmxWow6zkpK03WQ
JofbFLmO9zfJq660+HGuxQY6LyygbgHVAsao0pRZBh658w1wwcXn/n3NRGUTLoKJvtShxpyxhe1o
CkXflZ7xgNDSERB7DkUtMEZsNz67MwauLJrBebmYdg91c1WpJ4tDUCjGqfcZWdzSjkjl63iTQKXo
hVGrGZdjz7ZXNbT1b+6byaYIdbMJJCEsPZLG5bZoY8w0wrJ92TXIAkuH6//XDrVuHfnlbupfEbhn
g7sO7j0qcBjs/b7jsREDA4tMTBrpXe+T+5Jf2PrlvwfZ3IF++t5KF2RgQq3rR2v9t6tME4tH90rs
NM/sTs3c9Mk0bEGauy3PpQNR1/w28u8MOK0z62vBW+pLMp3/DVSXYxjHJXJI9ZVW7PMtv3p5MEsp
v76ExkyQGOA/7dv8oIGlgn2VW/M2+dnF+EauHpvuDLdRidZe8VJwoVl6KEVVYU2oIQjs0ynqZqOW
kZJr0o30E0AEai1nX/Og/SCf24OZjuvBQbXDIODO0d4mq7bOjXOFmkbGvYrfzyHP6zHlYvtj2q6Y
ODG1PaT0cer5jynwM+eIJXhMEfu2hgtY+nlH9BWL6jXMhJRleBcc6KLyjYxX00Y2AnMVnPLE3vps
gaqGffrT1P3IWKxzGt/0YpN1Y25JGi+gZynGq7qIG29S3DB/LSYQsRGAoY9zIkEPIJEaTwLS5vgL
NKmazqGz5dPKI7DSRHJBdixSROhr/fga7xm3vqi8Pnsz1f2/G0oJZh8SiuDskysRJWYeg6ZWQJHP
kqMGrsnKhalNZGQOnXMWFQ30hZsxlbLKWt+Y7bj70IEEIJ5dvG7blMEqRMc1uPeocgogeD2oqAWJ
BJz56A3zNQyKM3sK5uLgGtLR7hIUjLogJqD7mu1zdYKJm01wgJzziP625bpW2bExGhpM2B3eGRU6
3IbZnYN63/ytQEry8lVTR/jobOZWT6xUBcfDF75J8Zk8387jTH/DbDVGfZFVP2Xbz8p9xbIRZuDQ
TxUYGDHEIBf3wumaGHIwp77jyjUX5RnBoHGZW/0a8SaqNZlI3HDwuHfKs7i0ut/XfCu366CxpJX5
1Xu24/lpWf74B8YsLWJt5U6tQr3Xb2u91qPZUN1d9ieyuXLbL+jkDNMkkiV3o7TB/wg1YuwDqvtt
d+NX7OsgJ733Jxt10nQEHj/CjCQR1tqWtHZHaViPOk6oAhFHd9YWlV0LAezugBB8O7j9hbxQSdQ5
RJOLlqq2gFBos6CTmaASUYkje/F09xAsiPQOruh4dnLBSaaOOfWIN+as4RLPUAOc0jUEf/6a0Ul8
SPDtB3Rx9xoM7XAfyBMZiGHZnzvitO+l5uKsPOcmqOng9VaNuQmMTu+dBSh77Rh8uwMDw+wz0Akd
uLbY0jxrXoCl0pVc4e66vPaZMDciGwI0nuy5B/IdYcCoklsYAXiztRVyIPHpWWuyTrEslBKvTPXs
xEn/3dPP1cWVTTYxUaHOLsBWa9ROjpKhHh/7RdEV4myaECoIbruRbqqW10O3xAB9PFTMXOTU8HJA
nv4GrSGwK0880voK1Tct1GiJd3J3xL769AZlOlyasAIm3tizMCpc9b2h61xnglvlwrgDodPyQixc
PFRpm1g28NsLo5sDojhRnkMRDWM1BJZQ+gQF/yj7xfaBGUeUbma86IsohCu4RmcC4aqACM10BeBl
UzaWaBseky7MOKl6QH+H3zR7SLb4zYTeL00hCsMS2xJkM3flaGLM40E+k3sP1wwLfi/PYv4/j4CF
7kQu+kicsAgOx8gEtF8FEGJj5YiVy/dM59EKDE6YlJXFOZzdwz/R9Q/4W02phKggNRySjq6lpbON
yljHj9MBsCSAcPk4fpHEsNxaboaALqlYWkfEZXetHb7egUQAkqEHATPErs2JA3C85WoS1vPzXU0M
2pTwrRo5gkY85djUI7CJbn7YBMH/YDXgVOnLQnL/XZ915c0Fy8nWaF9JHjmwx0sO3Ug4nKgW6dTK
Wd77h46dWFrminnxyI8aNi9BOMWXqU6JsFjG1LWqeGvDj7HS7opRBS9RyDOYtaxaU1K89Y/B9cRF
SsmaFLx5n/J9187WVLIataphg2cGR7RpHXgf7bU8RgMgWWq2e3PkjNL2zLZwLe0ieJ/ofCgs4SUF
mHRtTf+rDtPF1rcO0hYpc0OBcrouT5PtO+m+keqT3XUFJukeOjDLPHqGC3i5/cyqymbxVHJBwWE+
FBIbJh2DOIIhna/4ldD3C0s2qNUX1hwbr0fO+xAGP03vR7ps5w9LLFfLsmbRJOdiPWdAMHKx+OGI
4O9JJ4q8JkOiSLHos8OxaDyCdlDMwOQHAsCa4LmYUvmcl5u7H9k8UhO8Lzdp6miZQ3t099iOLd4o
+IV9g4oS6FpuE0mKF64Mv0FOarj1ePi9V4JTeOIUXaucglro570wuhEcZDMb5GAuIE8hvLCaJ9T9
8RzGibDjQiLmjhZtpYrqJyDf5WtrZ/DfHz38KbvegsOr/ZxUqH9AHuTNQJRfeOx2305TzEZ3GKUP
8MRxxhzeETihDS2zvj5g4Uo2jTWOYjchmLTNZgwMhxySV7V58FQwXMAU1rRNaxlmUEheCRWrefCR
n9ZP2hoquCSj0qQeNbEdZPgYZbFHNtzLxqPiS5/VRYB/nJdRCbk6gBT7442p+145w/wgbaX1fYN2
SLcoFSq/auhkmDp2caLSMAclf2X0AYVS+pghdS550CD1GXOxfesK1/FLqx0+fx2qBBaGNWRijuyy
y7ZylI5KXVlqTK/D74f5FZDUxQoJSRp5gzLlHZ1FURemAGV0wgJk3QNgeuDBgqFyLpOfx8CFGIss
0s4oHXtlRdUl+xxkQjkCuyk6eVvILkaLejuikALAlDtGX96YzRD+jqKZGwiVJe3QYH1tVSs+D0Rh
Ct2x5Z/M96FKtqWcsBfdpSo15j0hl/jv6WAxFzPdpWabSkJGiBcN3vy1OY1e+ZkojuiafKAtcFUY
+EidJqN79kmkc0WCfIcHd2hRcUNjMJKbEIEIy2/wYCErj/zn+JczWckH6LbCGVauMjmkmAI4/Q+y
zFKJc/VQWToC5zyIg6qe9BRdrGOnLW9ojhTlyLPgC2BzhkCo1gPoB44ncdHtsBtNa3f3UDnoJh0e
FeA/VOT9pIOrLEYbXzOerkkBghH85W1CClHb2o4reUYQXi029mJGMXnSIqvkOA6FnAnmiDFh25Oa
fh2773qU7vjaFgGUzFKyX6XbsGv/1bWJaEHetRPqUSqP2vHaQy24O7tO+gLNXuo6TKVZeAmNrWA/
B+6dmyOYjwtwIkl8Wi9TFlMrSbyd/mq8mtm/pxDJIPeWb9hz7ji7ruW8H3z2VgKPHpfGZD5t7JrH
pG1GWZInsXPDlqwvY2NJkOvkfMEffaQICvqDYyMzEp/NJIEnkodIVm5sawzSDO+lq70POfw6xtgJ
0NHmmhJNRTlY6UlNmZr0AM+PnMEwJ/3prcCP004vEM2IK3/h+7fykcx1c3QCZTVeFYQdtZVA84Ok
5vwUVguo0bDag1++wVcG40WeVetSbUl2nmEF00txCpqnsnom2wK6S8mmD3RTm35+FPMuPrnSuoP+
wLPqx37nRcY90gd7CMRlTmFXXIuVc4PxoPeNhmOMpwi3W0o7iHRH34+1cg3SiKlxmXjgLs0fUav6
JeSpLiswhb0GnI+1M3rsAniwUTIftCtGHFzMdUeDC3qMQp+rWIElme8GM0YTX12FYBnmSO6nRsj4
VGzXTMYlOSP+CeppeTcSiBmcSU8fddyVIJDt6IbsDp9oLBJXAtdJW+t2jVV27a06SNANCeRcMy02
yFDbGdL0d/BbHtLXnevKJnykNpGyuRs2sNN7v4C1QEOb7JMFtsxb9wckzt1hFHfTIfXE1He6SbGc
FiV+GZRnWA7ud/ig2DZhw3pdGMJtMY/y8h9Gg/v4nE5cfier6bS/DoR8GXr2Y4+aM6o2OQmtu+HE
2FFFxs8C8BabCS0RvGuS5mRpjsLmh7VRf7etZN6RdE4hyDmn0yQ4mm8k2gi29TY1dQzlTzQlklbB
dAvYZ10SSbDBo3OVXhvI+ihEbygWc3+zISvodQM9kp9jIWX15LPJiO0sgUwtx7uxBn5TasK4700n
pjF/hwew7XaSifkf8JXsyGanp5XnADixvjXdZ2IcPetzFy5dpcqHn48szqqHhhAXngAycsqCMJlS
N+VtEk7zlavu+G7lkbZ5Op2snKvbB0d3NltnLcJ4K3Reuc46UTgg4DfRaxLaUyRyU5S6soRrF4Q9
Fnow8oauo5bigTBFHSWsM4aC1Tbwh1FSfm8bEswa/CI4mnyZrPL2eZkm7S795eocWJBLRDWFEhQ7
4d7dqXEundqd+SNVnGgethdoH+lJMJyfRnZl+YD6uSIUr/jdvypjtC6HkmXBw5UtTHYnQyMUgVeW
zvGN/q/76olBfk1cDBVeIvu5IddxOATn+rEp6NjUkr3eQM5R66CG7CApf6E/LDObVBcQunD3sU2n
ngt9hL2kKLvQSh3/JEy9X25k/TbhGorw8iaszBbpZWgDa3G1g+XmMbZ9JeY9g5W13F1AHYzg9A+J
QBTMQrLvs1WUKGspQVowL1G0PBAbtLgFZWpYtThbtJAWcWvrnOzF8kVIH+K3UyKM50qAe6kILZAn
KhwR5JQhtymxHX9NzgW37OcuVlWXgT/SQCctneeuLSBkAtM8eUEpQmlnGBsb2Z9ea6OwvJTLkHRJ
L+vbyfGSt3exT/VhI0URgpaNbGD1iNhvXyX4vr4AoWBdCzUt9oS0vkmQjVf0AWWcUSs+t9D+M5sU
NtDzeNXRotTl4925voHbFMTNhGQKqoQjsy3Ambk1VMk1AbHJClraHMI/XS0eG1DqZS1iLv8DjX5h
KJRIJO7GCBXILiXHqRcr/y5ZiHAVAH9nzF0zv61RliyA+QnnpHO4exTd2aNnkBWwzTz5m5Wi9YS9
wFZbDNWW27gJj3FxCErfB+vbqAo4Id7KKQIIk6FhBcTJ9BYzLsOCmNW5cK1dqJ1gw8E+GUVO+Mvy
evmmWbv2XVyrDprjuSJWWA3PeahGkBXUc4JU9D8KFeHDt+2c8q/YfGQ1pNxVKxDBNxur9zzHRBqz
geQ3cSREte4UGgzgltjhx85+bAbKbfTF5eSrm0VVVikmAp3v+evGO/ooJbaFd982AlrQdoz65nRo
GPYzc9PIyvWkHiOQMFbZKs+XVAuuo+hz2PQiewdjIp54xrx7JsXUry6D3Mdgq5ozBNkTsWSlORPx
1kLDjUgZdzhyxsu6lwjSztaQcHTar/8wZPdL+vnGPbhP8jPziA1ajsz/TuMzAMJNSc8cI31egSXS
96ZBPElMjKI9WaVXRIl3S+ETJprdNoPeg8wkdWPOAW5kbJ32iGUPEuJZzIiDGxIVT68/dBZddqBv
PbNCsGPKQFdLKDKU0Sd+9jH6ji1tSVD7S+wPmneSabUYlgPdqySh4d9GBkZ9p2suOPqDWR/aojWB
BBL+/UpXlq2ug3pM6aSJPpbcpYv+3d4TNAKif9nEfnJRYLfn1Qj4yPfKPwIiAyeejg89qrbpqz5u
O5mQgdymUNHUAw14ChqYM+zZEkYlW99nQIGUL1az55BVoWp594al56A+xqbv4VWa7T6KMslPft9w
b8yfB9/Xbm26RkB6jDSe3/2Vjk4C0vsJ2n22y93+Xda0hnNX90vnKJgNzskRzAlNmb8beepsNvPI
bYlkchdgNlXv1gAwys1vBbiFFjj6FUCb3dGKQPlMF9YZ4OUIKSHW8WV0N6MlCdAPsfiyRmDuB+29
/mYMmbLaB9XVU6yTWHo7VtFzGktTDEJjTz2z/VJmAXFUZ9dROvlc144i+UumBDNOMnHJpIllUG1P
Ymti5SSOCqK3z8fu3Wzw/466YuAOQgiWzU3Lm7aY4sAorKiXunUdldVB81N00owbrlyuTxVJbFAa
lB+bK3ZApkX7+g0J6a+nAvAioYtVcIQHtvdJdp4XS5veWwtihkic8vSe2siYS9WbSuH+dT5Gx0XR
hsTJgAuAE9De46mpWe07dhgbwIu7EYo2hMmotmX/ZRLcjv74tVlz02Ccr1gSoMFdjfCrlXwK5hHx
R3oPI82C4dhXGBcgBkeX0p7MTdZ9hH7qRgGi6aqHE7E1L+bPj97nX3ugikEyB2bufd4EH3HRP+Ye
fms4ungMdiczLGsgbcqN+Sa8MFRalJ234C7k066OaMHUCP6ZqzR2p90hvmSWViJRcqnM9kELI2w3
XE98/7NLuuuI7DWDdfJ8bEiLn/doC6N4w1U/NLLfGrn2rmT78Zyl4RFDc2dyKzgZtkPnbg8AjScL
A+1Bb2+gK2D7zlXW36h0h5ynWE1wZkwXjUJfEuimr7M+PHGUXSiKeq4QtKO13sNxmXgeeg90tf1s
3eHfWzVRJm4u3J14ZkgixE4Sdb639BB/yZ5+GJ8q3TRdXYP7uryGFgv299g37dQWrPi4EjEG5unr
xh36biOzCq0LFxTs8ed5cHO0KJ0/QCHEe6Ev+7b9ix4F45XOx3p8DM3PVvOgbG8XhVKSv0VA0S9T
YWuc1ZUbeJuHsoyZdhyk0LvTuTNNxYXtzF5J7Yt2ibBeEkVtQLy4yISfUekoWh1qdDcQIGMYFw7r
z4iHi9bLOvzPFwg/GU0CJpiRFidAbG8UoDHWxQ4o/DFcQMGqpjyaJGJNdjt5nV/UWnP/rQvbnioG
tp8Xp/gnt9sCqDce1d1f2dxt2kDKT2Kc52vjaeLpKK2Te3nZSAav4q6fZ2600HHnJbQqJvU5KsTU
yNu71KEPCSs9dp9B4rPeJOVOElO+KXU/gWxfGKPbxcol5V3NE5XNWcAHdCJ8kHkzHdERw6Y/kc6E
UjQkV8pBaD5cyBT0s0KTw3WwLeVNMAaMTQKRPDnXUrq/lnid4kTtpMx0nKAr5twPVp8M0z03RVfB
wRpWtmytkn3HYdGykSBL8wivTNw+hxZko+UJIOl8IavS9SSFd5DONOygIkDtwtm/KahQTcZg2TfR
m85j9qIpOyqksRta5Vuk8wJ0gqvs69wa0YPzB1AD038qHd/9p6yH7t/Da25wMG6OJJgADBvdULPM
5l77sdmeIzgXSzZ0wnbaP78r26sINpSpGPNBEGTnvPLolVCP5v7c2KUDrqlQ0HceSplQ6R5ZhZKn
tbcuT+GL9VKwPnMl6Iob0O+kzbn55H3ecXPqFbs4qp5JTkMjklhG60HKIDJR7jd0M592lgCMsubm
Fi8SHqfXFQLNP7NhS3k4L4IKh8te/MvIUe/lbomu1QsINfZbF305TO2378dOJipz3kBeYZrjKqaE
Uqda7BgI2FMVlnYTVyInU/oEfKnZBpb4cs6Te2q1sfPEVKgtWqjmEQBNRkQcnRKCrRDjhvv0Bfko
d5n4Ws9c2KmlvIyY1b+CZ0tJfUcJbuXPpAX1KY7MMMVBOCnf8w1NZ6E1xS/DIqCzoBIrG6HA7WSa
V0KPGSKJyw/o+totUP92nQc0z2GBQmtZdebpmSy1PD+uaJBmVzQNYz2sMPTqGtgKQeUzyiFCZFFl
WtMHpO5DywpKmQ9ROwQZMylLbJeUIAXJpfXzk4o9Ts31y4+0zJvwPie9oaQZmxMs6f9GHE8bIzeK
dVHJKaNRl7KidZ54aaURxoa38+uygTvyaeQMRd5gl4Zffgc6D1UQOrRPwoFfkf4tAbBLB7p7wJgy
M+hamwBK7BHGIjI07Ynq0gBEljjtLoFMag9KhchQ+Zrhu96nnIf5W8Ml9OWAtUkQ38IMxwiTLgYb
N2TzZBN9ljxpEvvn2gFFZmHc6fAoUob31ilxq1P5IyeWaIH7f1SLFUgscku8bxjcpronQgdYYoN5
oSH+B5gZzQWkmzx0QY5HjB5o4PylllXmhVb1IQC4hSyMduLwCR/BqLfTeTMjk99Qmf4wvnhUulAQ
AZXsWSJKz7s69qC7VXUO0/F7Br0TuwPUzjfbtzQnh0fa2PgjNY51ONasW56dkpeHy4jAAC2DhQ7F
oBtkoMJSDsGetpT9+YgcqOLTqRcshkNA4MLg16B/gFRQu7UCY6Ul5RNbGkoz7rVzfnzfIX8ZYN3S
cBeir8OMiudPAomT0gFCE3tk2LCmZ27gEVx5rKDA7/oCCHTcWTCIXPu+nplcH2HHihO+pp70mHR9
5O9vvDbLl3HOL+4g6UsRxXoBstc/VNhuSY7Rzuy+sUzMygQIgKbwpQfPo9uaiMA52JNZZxQ/hyps
AGhdoA1M8rZ9jmwOgXWut9/QP3bFW6wo4iQl7BJ2mL86hM9uIDIwDymhd1E1U13Kd2Q/D7UE8s5K
3gZUTq0KIDongHJyd9ZRKg7AhbkJ5uEu3+ajkWpifjGJQ1uISyISAKXfAqSjSO3Y+f2cyMkjJvZv
MPDUTW1uebUJ3o5/T7QqYxRwiMcAmPGOqVoRsKLnoEkhuM/qHtN6RvwV4zmMEtr+pC4KkIPvegBt
0Tv2K+9O+tVJD/t53LxC8kxbg52h34ju06avri8AQaiS/DF/KxBZhQH0nO2eqx60zfVIcmVA5tNt
ni8g0waNpwwbWaFD1dgda/5q1olnCFLvgmkiwSzV0Y0e35OaAZW6v5LtAXMZdzUiQj5UvbcRqMLO
DUzaNk2i0RM2ItxqbmBrqnwTyxZh6cMWtU7PkfKgjoVEAuuacl/u5lCjgyF4JnU4BTxwDPK4qCD5
V2RHXGiapyteowoEXDjvoMeZ77s1uncqVHk60ckb5V9ruVpVxXO2vR9T/U3Wsv4/yELu1qyT4qNo
w5IN1okGlVY5LNdqBPuqLa2lNdpaJN71liFeVJUiqAeM7ZjbobK0ZoR2mFtQqJupEUv3y0Fjj4sa
aDFk3T+W6M+Nv6BHL3wngKlGkobRl1TnmStlLEkYq/KP/sRmuiVAMz0mgv2PA54tRO6Oncap/0YC
F1bIfQrwcjuZo+kJFbYs3jfpUQtPgeKTDgto1QuXgeIJcVj7uIcDwxHBqYMPmRAP2XQe5OBv2NHp
Xv5kCS9YwiE0zix89Vn1l9UKLxsJEEv5IBro9Tcx7b2OYM2TQLIfWV1CkGUkfHaAimyvGG+0BNY4
XS8AJS3fn7T1lXMIbsGjTgJSI01KVgMh4Uf4J9PLeuRhda6gXiZDm8Nn1KkBAkZIWIpzOFaB1KFS
JerUO1QP9iB9uWKaIkQ5myDqjH+LNFSNZIzTiAjBuPSdP1NoySqmOfdT2q2u/q1zQ+5TtNhoz0IE
hWAFRBPyR6A+zVIknOyOAgAuWw4e3Q3oqKel3GwgIOrGdez8XdkRE3ss8tXnQKusZNsQc3APUNAq
nbANqlRJMy5rAhAgT9Oa7pBTtjd1PU1sPlG8svBKO0aCWZveVsOZSRfV0fKA5zRDkdzMDRkTMdDI
Hq853c2EAaTNnOn5fKL0Pay4959Tka1sMo5JSqdydIMbu7ZWDBJldw42uZECqhumOa8Di+wMhah7
jcZPM8F2eOJVprLb0QlnjsfnKnDz16BaVaAVJ8KcVTxQqmlGJGsmFamEhz33LszBev0Y+QUNsh51
FBIyiJkL8O6jMu6kW2EoPoDSzLoN2HYxRcMzcyDNIq0rooZdOtgGjIfNBpVoihBCx9OtqiHkd23Y
E8vFK9vjnOu5JU3zUHNRTGDDh4i5l6A3Vrt2+IxHDqHJ5/2ccU3zK7ihc2Yskn15u2mK+1USpRvK
EJAB9h1dfMKvIy0434sdOHQc6EZQkLm38Wd6vYIEgCNnyy115ZYHbg/A4EG3izxFhNL6RxIYwBzO
OPZdebbtmJmgGvVvz5hHnYnNrhmthFfZedfQkIhM2XS9uaMHbwsjtaASEIjYrflnf1vRJ/4u8NRS
A5lCMKNvKpwNddyGacHVMxs1egsZEpnly8KShYFbPfR+cgunLaOBXs0XK/Iq+R1UOQpMh2piQqHX
gE0kITRHRyXpAt7XxJnH6jwpPDiGyzvS0RZFjgNW+01kckMZNDypE4LeCJSrapcCB0JMiJoiFiNI
Lc4d3AMtzn1QmzQ5TSE63cahiE7hddOKN3OiN2zNlenaDBUrR1m5YkYCvwaM4EELABFwfuA9DNPu
O336Sz4YC5sCoGO8hjPG96pJbblRbVi3tGkJqLtZXBUVJis2AwMioLW3u34LznPdrwEIOIjVnyfF
8eXhUnIvmfVeuf5vbbnmmJb4dakzct0rOBjNz9qRo56pdhXWidLQIpXBvr7LNQHlDspk9kq4MwGU
I1O/uEnf+iRCB09R/xNammptGHWmunFy7VFK9uGP2LxW/QVKGZ0g4uj+SLAhToq6FhmHT+QUU4ea
Is74La9Izgl82DLUfFs8m/Vj3++g2T1Jf2kr/MAAoARLwWRzngpubMLbU+p+AJESvOVEZwzCBQpE
xePAP+o1dDQBvrCrXULghrOVnHFyVf0WPMwtF8lpPaX405p0qRE/aawpPeEFvR7c5H4RsLZ2Pq6s
bG6BT45NE2q51Mf1u5MWKes2fZ7sLiafToAkDxgyn3HTZ8oz4Ms948+6okhl64yv1Rfkdss2yXqU
peyJqM1Mfyvzl3HH+8uniecQz8fv7Mn1T9EkN2ENXF/IU0p+T82dlcBonhiJJzzV/ug3rDcc2CGo
aUS4PJ74JoJTTreJ/9mlR9HO2TjF5R3BgxTwdho5sF+oLQ7DK8KzM53PptFHjTb4TcgPKowl1HKK
fSTzQke/rqkFgVHKFyOGF+Euxgsel5VEh3M+GD3cn0zZLQJr4Ljug86Gq+JPSInIa5McZa3ljaTI
tMttLUY8rV8HP3HeG60rd7zXYN5PdGMs6OGKZHQUR5f8CUtAR/wukcOJFh1Jmes9w2ql+SM/FanO
JVtaHgz0ooKCliKxEtYgRdTA9Jf+rYRqXRRbEz27TM4ytVk6rGumU1INvk22dG0fIPfk2WeNAdDv
In1bBxA6dmCO9E2nsOyCORH7Rzz5deyAmBCgH0MpxkNoVHz78byiuoxBj4eFzTfgeDYO/caOhj22
2pxqmt4Xcy5y3NZGp26cIEaDsHyOcytVXZlAaolqUu9an5mUK5mhJHJmlcyKtCT3nr5QSSMTgR7w
7IXnABeyJjJXnYR3hT2vBBVdum4Pb5xmypnDVB+MtXgp9FoxPUmOhp1Qg+qCEKo1NLKxAy1wHCfg
6zQq5x2GDJo2h/QDLYhOF8VI1bPWHyTNN+n02HImER8LSUUm0n6Zm6G89ndcFqPXcpPWd2I/05c6
nivGqHRTEelJeGPM9X3Z8nlk++06QwWiJyuNRabiJXC308i7meGlBMPO5E1Si2GWiRp5WJ5AxgzA
Qiofy4dpDq8DWHJmRZozBtAAaBCReAQM0RLGrbTHArp1jKsVN+/w8fg9S1A3PrVYDiXWuoogojh+
1coxEFKqkAjbPLO6wrAHEmMkNZNSWHlHg7hGNeMqwtIuqIjzTX7Oy7txAoDht6jihXvvPokTwPju
Ls8kF8+88K4W2lwpTiulzKNUYOQQQCdn7G2898g3hgkIdoYZFqRrah6lNN1en8qQxy7ALjvQDMxt
ktibkySJQNhzlJGzhxRCzmX/Rir7EARBefn8+CATMCkBiA20lm/NTAQnp3IdsjjDGts6N53TQY2a
J3Qn+LGOAqORDRdadNWA2trRNnEC8td2c1tgBGS14kmEA8w/XS/CCghtZaXWgMne/WeMZdmSKAI/
Zf/b2g/EYP/dG1oUyeNpWIQl36CMFgG+ESae67HyrptySqMer+RK7Bdz8E/bwHWYOJKW5Fdv19DR
s/qjwSAGflDC6ytIAtHt1KFzYttR6R29larUdeX6T7HR1gBCMuC2aD9XPTATytrleS9b/VZvEzB3
gvHU66eAfeO91hxaiiRZ+zPzEHyi1Jc0sZ7WK/Hu8XpJ6dUTwBJNPZEgdxiOhalzeD9tcSBJShUQ
DMasetHHH1hfBmvqVdKVAObQBuG3p5Veh1nGuVUUG7I2AFmmv/fsZELH6pMn9kHbnA32V/x5299d
kMamZKoOtY9AS4mreD6iGoVjM+GhiWcttJvBaNjxYquvJQTgSfozitO6iMW4G6Eui/mHdAGS33VW
BYWIkPDzSZj1XzEqFKVaMgl3YYI5aL0bHq1WQ0i4X4U4l4ASBWlr8CfnyGD2AoBIK9QmAYt6jdsk
Z+0yGzWNLb0K2VVY/Wt9HbEaDYg1zBdo3jGx283mX/Qx8qjCWRN6Xdvp30tBH5AXpdYhIfsdEHPg
bOn337nWcD1q19oXWkJMN7sHx92SaN4HsWR2UN/iFQhRw9PDiQgUryFON7zGJltmK0eRhZ3yHcOP
eETGx3OT1D9pLU6mbIWMkM87QBnOUIMsU6aTj8rVpk8f2+uFt/r9aw6R+uUlz78QFic2VNvSTp1+
OtwqY2PeG3KTRcTLhKPzeKA9qtmOsVkw8uuiBCD+Wrd45HPfaVNRtunJtjMSbONM3XO1iBEZzr08
JRW+3b0RYNmssK6Y3JgugG9e6QsbwbaaVUghou+3YJFWWTrN85nPb3h9srseFHtgolF9G6t7G7BK
j1hIik3bZS2+3gk6b2ZDN8A1XvnZeYcCxyZoQpavbalzYOqGvyv7fhuORMoLel7Uge3et9Mf2hJr
Vh4EZSDi/5Y6GBOgCRQ2MDVzmKAF4U7yyIle/T4eTW5cNVwndCvr7JZahYcmDelZt6GLHkaS1aaT
EbEdMpFnAlxFk9UhwdWRkG+ZF7pVjYx0oHOxpI2hE55WWYEGIzoNXUsr25q0LQAMi90KsG0fTGIp
O6ckqaIkGp7C70lAEcdemGc1O677K2EmBGlzTJlSzso/EcEuRRvaTYxj2hCtGSRCIu8EMDeqIe6Q
NWnL0r2ABoYw7WloFtHjNqdjaqKO50HYcxOrWWwx1pa28b5CPc5/asd7RL6Ed0KEqD8ktUcRcyFW
o6So86NPZZPbWXZcnOXQ0P7FE8tX4T/nZxhrcDw397+iWYsdpO3dFG3uQDuOb0okB4t8Q8VXpCsO
FN/fhm0/mRFsZhf5JO4yRFARcFt0iaXzjKgRCdMBt4xzsO7YV/FG9+bN2Y/sz/fgo6xlWjqc7eXK
i/zxfIpA3cBsHKNedbpse7MSltxhUjyb2TdtfeiGXpZRgmOgMKmsxz9mSfMwCPcGDTjexdRaahHu
dwrk3N1RKVBlUeFBk6LJ/AUVcZ1YrxHAq8Ppe+aUqoDIBPHRScW562Wr855wFlTk482Za/3aF6JY
1buE9UlxZmWUxiLkB4abG89qCgHS1A1D6WLpI78s+Hj7VFF+S+k9Tj+Z5yBmJRl/DZfV6lq7zBeN
cVqbtK+Kj9z16wd3KbpYGsuI8JjfYvKTna+PN5xQLFVdMcH3T9wMBlfv2ezgMvT6gUWwDPLV6/iR
r0ONZ3FpTdiCXf7rQdhUyn+kj4UwHky81lfB5LcgdsWojWvl654qnhXjJyRiHI2hRcXhwnPLHwW1
XfYC3O2NEOZa2se5zLKCw68Au23TiTm0vVCa3VuG1rKubkgmAJSxGFjn8+Gi0RC+fMMFFF+FSLZN
VOboZQbJehPW+ZhhndDzzNnq92dkABgYkpK6HRew6YRnNXshsUpWKLz+35e7ok7n88KU6k2xtpaC
BNqqdnBsGiJ6rixpTkiuQFtWS38vJzQr2XacrNA3h9gOGMRRaNvBBinUwgB3SUe4XUVoJ4nnsM9X
0vg91Ufbj+aY4A8B41DfBSFGX7pMbHOmI0Q8zTz5ftWf9uPJ2TlKI9UOkIESkXKryc5OKvenX07h
ageHAeuq7Cm2tso8zqyNpzU4VRMWtIsC2O8yreu2rGFBfonfkxyLpC7UeQ5/6V6CDBetpbQGKzH/
2eYxibC0a5SverXXykCzxVQRKtm4A6O2ygnVeun8GloFCHR3ZzX2+gZybVOy5VlM9esPaqKkGA4I
ukZr2ZR3t0fzKRfiL46H8Zuyd8bAX0lGI6ZyLjjoZQbb+ipAK5QTjaIBJCzS+N52KCpIIT0IeRjh
CR+BGWxYdPtZwUUMTdwoNW6tuWX91OVMgC0INqC7EIqrQ5jWiWxisxbBuzUagHQZSQwRZ5VivoOo
dgLKus4btN9M8Mol6dEVlflwWcO5rdkeR+mzsq2DesKPPBlSy4gwrVvIYUYt65sKdQ46obwSbXT9
TK/PzSXdFnLyK6Sw+x7S1hLri57W8WBP5IXUk6T5j5zq9S0j6qgPurn2SIJH7PiCox2u7HaXAboD
SI2RIu28U2UutKljetiqjkwwQ/bFmI0/lY8uq4LKJYeOGhJ7HiwdWtZ1AWeBHsTGtCqM8sDRizql
CYfUd+pqVGSwGlzf844kAsG1pRR4IMKbHr44XaBuOtVKcDvHl6y5nG/WMimY0P8ZXnuQ5qb4diZD
T0qTJ0OFuvbmp8SUM9etVTvueCzbTSsiyth+4eq0j1Ofahm26J2nfsl/tcTF5Hp9Czq3bw90bFon
Fegv6/yijYZeH6sn8VndTtoPM8Kq910vWeET7Ni76Oo1nazCx+tGT6c51ecI0LY2ZZWa0fSPxwC+
YT8CitEM1EXI0WguVUqssPuG8oKPnBmJAklKv9Vnena/7au6MO9n+vRSKt7vOvWX4XQF8RB0QXGN
LezWpdgV5FKmZ45gQKWxumnY5Vok5/t2ri99nvujkYP76ufqkMoZdA/I2ZmgE/qzUGnEVG0FzKbB
MFQAt/NLD2rHtNpshIwqIdtFg7WasEYaigJYSc/9a3yWfDJ4JrVkWstWAEk0iieO5rGMf1RYIV96
YMpemcq4yg7lAv48i9gTMRkCR0QQrnTw1gp0txppl4LPUa5nSUrpGgfdC9YgGmuEZrMqXhXrtO21
6wdkTtokX5nW63JA2VTH5OmdbBbroCnJ/ufQ7WtUOKdPlZa5ndu74EVy+GMU7Xqyrnu5zGg5r/h8
Y1gu7NQl4R8+GPOCgIqD8dDeeA/XzmxWTtHOqQgFPLgpPlTzFoipmHUQ6Jvn0rbdV6DBZGCMTIHJ
RcAolnEsvl/XXyTcOz4EVgF9LbMBXL1+SqYk+aP/o1Wmof8T9iOklZzZNsYNd7Ze74nfE+FrmVPz
LatTAubvu8neZ3USK4FAyA7RII28JFlMhfasNitqEGyB6IpxuD0xX2Rd8A5W42k/rZj4O8d0gthR
o+lDK9ceMb/PWr0oYEp8tv7/XvssamJTCuZP2SwUtmb+V02XGZmMoVzXn75XCdi+dvO//90YpyqU
VI1KBPj2mIsq5shHIoX3sCOa6W6wLJNq5WArBGExFXQVk1hhiCAdYj00+MQoABG09stsH/m83OOO
mbFk/At9sqhx6sh5jcf6Vs8Clplb8rMN4txqb90coY4SpkUm7w7WTBySi4QLswlO1h4dlD0qxHYv
+tjmpvEHqx03tRCpVJ+XTdCHgOwmWdjPeutOels8gNW/zruFOBQRMmwGeV2swRZNWTzZuSdxuxUc
ahlWHyFcctj/KlUOvCttgkntSWvf0f55WQ72xl83RCbH845emVhXUBShJz32EuZir1fAOHfvU5f7
iQxiNIWQuVy7GmJayJmqd5sCtCpYwlUdkeluZG6JgWm2jDpcCb4A6Bp5KxgpWxvAaiQ/NjgGEMV4
cdqy9A6OyyiGQoIuQ9eNNwz9Aq83/WLbuvO9TB4PuSSoJSqTRx1wpUvMbcC76uVSDgfYii/76HyO
yBRs7kNkZ7/e4CDnrcZ2as8SdSwXdJJU3FsHvmc7CrXyJa6htahplksoTS0OSWMwecK7mdxX6cYx
2Ea9MhfRThK5lfs3wBtQvexRAIa/CP+yjyaz6Jb2WYFYtdmIWw+ZAr2+W+fOX8sgFdDp1b+tPEUW
0sfX2SiYIZurEQMEhBk4I8B2Uds3fIVUUaySkqeKzC5UdM9XcYYNzp1fgsCNk86Imfth8IzdIL2J
MX06vKwyBK1hNZSI/cyPieqxZ1qsKSZYzieIaQ2kbEsiZAUxOTCjXhAbdH3T2C908AbctSQouTEN
9Efv0BbdPZt2rBDsBAx1tciaQWLsMlWrrswwB83NPGT4HQ6mdJ/j3/GH7GpX3RisMN59Svbo0klk
FmuHF71oZAHy9oq1/scnU+9Z2G166G1T11+CbAfClNgkzf1fDXyI/QY1FMyDYig8/rz40SD05OzP
59M4j77EKCqDOO38fhJpp5VJXicE08D/d7Lsvn+ars0GBUjykHWlPZDv3+OZBje+egYsdH/aK+E+
cf8sUG1j0JMHC2kNvF+Fh6N8/Y7gG/cQb77vYxG+0JhgiyyDL8qI2a7Kg8/gVwr1bJlozegTBziq
lHTxX1DA29fwZ9407Jklh0stcD8xPnumrTDe81zX05J58ru6rXGfydl42ugY2gNENPeOaMnnGiVp
5FhiVStlIcrLm2YlfKDjcyuf72XGtVdKSX0ssNloKsDAJdzguUymr3uAlX/HEoWDCcRIyC9jtwxI
cjyAKUkrcXxrgk1Qx+7DFez39K+lDbq9hOyRGMkE7UMa6LSDGl0tTAjp+oDhfEBHE9yJF3BG6z/E
Idm9UffZGJWvODQF15MDt9TKsuvvKxVg2yELywrFSZggdJiwtBKootkJuOd2aX2ikBRGopxdmg2t
dVWm5w00Gr1l7LxZA46RaOvXuPyKWWLvefCX+yOiJeCX7Fxdv+/AQRm6bY8q/Lw8c/2oo19tjIbw
mDDRDte0WyOzTFuciK3mjWadJ2IotpixZxsfPHHE9+N94aOR2D2EakhhpwHNbyrzyhPonRQjTEBp
4Pyqfyfdy7raPKbBa8RYEgmZoa2kAa9GhSJOcvQK+P2iNVJsZ4tzP/KlT8F+BwAjC9NLZA5CFb0o
E5oGJFe+rp6/n/YS9cs91elpH9kmzfa/DtTkUdTL1k9rTXCQ4J70VAgJlUqve2e2p6rxzN4pP/Ua
O4v0jZlJ2EnAjxJj68ehwOsQw2Xu00NdIaHvIAnFWepHxpnN1VgZWkmhAUOwggzASmtwrRtEXqKN
OOd5kidqGDeV8afz1H0uskCEOArYTr4R+oQOwgEgo2O7IVm4VBJ7owhrNUbdrhYgfzmJXy0uIYwa
YjuTTwQfJnfMzQ6lXcdZKD4QzP68PLgSa1i1K7qEJ3/DG5DzKV/s+bordRfsjKK2xCmLcCp8jXEZ
5FysYGePsh19Y7UvAz9AB/al7quNyRhDXUGwSaDe20BovjJrATMx29u2hY7uAFLoA9Y3+6qKCJZ3
D4Y+Z2VhxQLdsdKluQ6SgxZn+4di4aUKQoHWU1Vng5Ti/2DfRV7EEmy3VW5T21v/wzKVcfgsmUIs
zkYkdJORC7cwJ5yHC+07RQmkW+wMz1CXZEbktozoh3n1Ko1+GwhU3b+Uq6y8ExbCmF+DwH0pE0hw
ywHcTVF2HIZcZPje/CJH9CejajQZDXaX6PS1TDjJW0a5JVmCrFTLN2TYk1vywTzKwhQte3NFmYkJ
8aEldnpiKsifNkLPPMab8Xkn1ENSdlTkN43Tii+CmnUyMRBjG/16mDkR5NXKVHsx31yqhW1U7obP
gOF9Rnstafl9r+rjS6Ym32Lt9/6tYqR0FlmXeHq1hCaFF0C96CqewPWelFY8/nlFAUr27QHfHeHu
cJF5/PsYlsVdxpG3AGC7jpBYyW8aB/wdrZm0A5UuLxxRTi59Kfdj/+vdsBGwyAS1PoM68/uvPZo9
bJn9wUX8WJ1I1J9z+4O71bo0iCF/U7zhadpMEjtuP3SRMa8fOtR/lBmWTDbbUURBWrM/Waeo3tNn
KeQ/JnFT/5jaEC3Vw0Skqz4lu5YyLvqED6bLjluOg+GKZ30jkAItAueteTalPtUzkkXkvoqFLN6o
TdQbQmtEEeH9eM+I7CzgGegPeuwqeQ2QNnwq1q/jyQnKc8fDdvXZvJAwVx/mlmEl1p9M6a/ZJjF2
WNVHAUCGFmny2U1SfspRMY072dul3l4GLn6zOsGwzHJkdYL+VCC9kbD4FR2QngNbvw/c8tbRN0UY
bUC5/VD4IWJZh0mNExXn7bNhBQwxLnNvxFfzs0mefqg8S1uKPpsL7m1s2up8VNpdNapR8GUyD/C6
LfjtqnoluEv2QNiFHc0zsyLD9vEAa2wbqGKum/hAWMdxMz4P4IV4C6S3EDFRF+7bhPdUlGEZrIZ9
rwEC4RK7rQQw3li9aat6bC6nQKzska82y59bLa2+3ShD5MdaQH04l8cpeGgU0rXAlvtGOPUnC0yP
gOUAONGbR4TOD7hpkoXX2sRtgDqNvm6IGqYrMhBv+eNEFmvIeY/t6WDW2ZNDb7pWWDkl7/2kiuEr
6+qVHILLy6v2twMVFy3u5i+4SudNs/m+Nzj3n2khcvV2+dbAqXpipM4i2zcX5AvFuowEPL+DJca6
I8WhS46cBiyvmCiq1yRGSicFZz3CoV1gxn7XYpGOVYaCwyi6ZKlBc0KOSs5w7hzFsDas9DP8i295
hnVkqyS1hNKijJ/i0tTRRaGzvCsA8KvJpoj1BgAG4Gb+5JXLlw0xEeEIZ+kc6vpBZeeIkV+scC1x
cXLS1Ycrg8TXxahXEYt8FnVyhLC70K2GFQw6p9IIzfz2QWrU2/ffLyoKsw5Tl5hGaTJm8l3J8NOE
xSrVbtcko9VJlRmPwr9fF9D4ylKSu3zsSF/aQAakj0b5tWSLpFxoX/nNrcr+O0kJVXqnxvkBrJZW
LHNbT3t3T2HuXigh9lxNF3T/e1NSP/KTZu/kZVocGcTvC55YbOPAYECVThtKGOfkleAJxDIjBcSM
ayDae5lVoiKKnF2U1hIui3Tlt2JZpk5oAMMHNWLI05/AMkycP6MddqCEqqzc8qp0itBmoRv3AdGW
shgiYVHpuujHXmNwWfcg95pP+zuhPnpWiYluqfg0Ujyz+5+9I0jGMf21UU6rVFe2DpOwOX1inH3b
LrR9yBge+hDTAANbi0GxBBln0mJzmXYOmoV6I9XVE1UWjR+ba7C3XpewHOJs/U4aX3S2BBnbfcPb
VohZSVR7MwJs7u5neBKNZYcRHA0RBnpe7W6fVkF7OfaJOwf7iA0ffF52Epi8TSez7fXKGL5UU90o
fXeKXMo2X7x0IHcy6AEqGtDSFEnBUNFg91f5TwLkL9it57HHkHKy8EjCF4f3odDrAdwsv3bHFETa
oY1zwX/SCKc7cp9K8kFb3wh9Rd2xpI6i1nq6FdOnAFZIQQk3+u4ClmUgZXsFkjeDkAkPhtKKwmlf
42oGmz6Z0YtGVljyNmx+Tp1F1MBxmPdHbCO8XFb9riRVbb51nDr23vaEMifm0kCW+Z1mSmccwuOE
ofrL0RU8yfyrPHWquZTAkpQXDFEV9nzu+EJbnyWJPN9nWF2tbr1/Xh9+pq7TEYqhJhaBSiAaHevY
GzL6bTiHUBSeJbU8DFOishV8bSxZX6tqiCC+DnubNJWpONrL20vO2W4CdzCPzbMWRdNOwRf88vCn
eXPdG05e7tggfs8XaVbCuoLRTqAV0KOEX5+gABzW70HYpBZIrnLcLp9ootD9V2XSO4Xq3wriY8ZA
QuMNNn4X04QSWUoV/2s0mC8X6otBwox9lw2fYovWV8MZzBGG5xtdzMfBMHVPTWVgD7VcjHg4nNmk
qaPLD3SO4ZUK0b1jdh/9M1tzAmbiibRCNJZ4Vc+VZSu29vxeLd1vKBgWk3s2srr+SOmffcoPtBmq
m6ZnAxT7VGRkFpCC6F8zdFchF5mDF0R2Py3uz7KCm0ICDohzDp5GRqkF0Iq6a9RNUlEDt3xMV5tj
97Hr+WBp+BzAe/PxGi1oAVan/6NUW3bdKlfjtORyYGO86+TnpbCDo+0WdxR5NA9YcPQUJVBTQt+O
ZOc1w6iSdd2Mc4oh5gWR2WKo2bZalhL3qhvrP+vWHXPyR8yHSgGLgj+46fY7a7lZOtJt4C24hNup
+rmlfct3xG4dY+MIBBXtFdwqL/tDhFiEM3/DR3u5pZD56WRmF67blqKhfA8MjoqGb+u1hoFBAhJH
+IsWLZXkvd5/Q7q8kBiY0Urzxgjfw+qmVExX3izeRWAg+8bgA4nX54nyFcVfHbEy4Kn+7tQipzdT
q7hw29x89A1/krLLpDOfJYQOnO+d1egGiCOtJEcYXgkvnPn3buTUuKjpbp9BAinVMnuonc75FQJC
ypU7vqbhs57K6R9PuesptrrUh8oct8FF//5ihr/VgCgxTVpZLFdE0nqCZEn/dLzd25L78yxzO4Sz
7aG4ghfdLcVtITFT1dYuw/miLC5lcOa7Ly6FYpKKk+1pFwQ+YLvmvlk0/6QVvyNG5ixsHpgzGtZu
kjA60jqSlik0a5F9hql2iQGsYaVGXTQzLinEgCmhglu1wJLfeCnsifZJp7nNP1FWOESrct2MqqcA
ddXRaSi9+SrOQIqtSfE+FlWrrW/EcPxu8g/zaDYBQqDh8YH1VjvCUZRPKi0sStHOKmDdfpaZUoQw
xzRuy+cqt/uggAHK+WKFWfVgXyP2a+AoeeEqlSuQN2JL8kaeyHtkjg4GA491NPWtg0Z9kxUGO0nv
E1yTfdUcnnF5IoUoYCvEZd9/Bmem7GGn40yY1SZ9KXbaC+ohPPzo/835tTmS/rE7V8QApGx35qWH
TZYad8nOjTjY8bem0yU8vBCqlIylzTSAA/BmVciAaEIQEE+GJ+FDLDUCv1Je1IJ1LI9GBTVaIPXb
AXeiCTvXt2oO5/IGq0bFrOhUdUvD5MXb5j/dcjnwP4s3guFuLPraWTKCU/meGpGEUrioiB7FVWGu
RzArSiUhQVd1pAVZ2jb5Szgzs2gAnjQhmxK9qKru5/XSMi5PicCVcGFyioieWE2JKU87ICBz7OKQ
W0qg1THDBrDIU3bI82tIE6+sh9h6I8pNXtGU33jHFX5Wmosx3RMtLrKPDHXf/OXyuHphNmfqR2a1
/eUxtebOvSw4wiThEeNEIDTrw+pCxO3JGibPgRE+sAjNFV6cET51hH2+tFWvrxSN1FN1h66M7Q06
xXuieTdApNjky1VIaBlXsegDcJwUuzr2grJDA1ydNGUR/5OG68P6WLcaS90ZLADBKilC3w+AN5vf
lW7EhxQTw9IJ+PcJvd9aIqpTyxYG3SihCordoeY1p4ypKY1f+gOEzHSDwwfD+uiHpgfWKzCYr5xS
yBlsNVYcrTjfHo+w8/eZibM3KSg776eZObaPsptbMAAllncG5zaRac97gC9DS9cBCjP80ChsMpEM
uP/ME8UJQMP9v1T5GE3Qnq2Iij4Ayly8TdBsba30/CPHwKTiWbDE1EaSwWcN679NpiAdMZ4W0nZq
HLQKJapwxYQwZwLEHsbj67lq2saW+0teOIAJLKASMznCGNZXfpgFXJnffjIKA/7oiP4Tlik1cAEv
XxK2pJZX2QkI7ves/QUb1uASxvfW2NQAtvfec4OwTDP2UlBovHQq+/Q5dAIWDyD3bWdRa9pH3XSZ
VtMhbpfdMfbDU3qDXCgEh2uNFTarYrTudYUQyU+O277LHA+GxV7rDBZbhP2zmEJiOkkInJKsfW9U
6rekg7av86fHBvVGubPVUtNGOg2U6NF5qBHBHRr5rFtTPybqtfaZq0GV4OaZGBIAS1m9z90auiyv
QxufGU9i7eCL62inCS3GCyy7jM1ppA77FlwR9SrcmreBP9VEUOn5qG7MxkE9K2iht6rBKv9weAXx
oCEzoMko7AJfSz4l2nmezot1W/duZEgD911TB2tLgE/AOpZNTp1FYpp4/Z6LLhAl3p4je4zkU47u
ANCSoWJ28lEqmSuKII4+I0sSmoGtreXavQfIvw1ZjRU2mbpoWGvUltDfjPjWrw7Gul7ngDUOrx6a
e5z/rQK8Gd/Pji12nSYf/1NeN/vAIR2Rua8IlkGgfONJLC91Uc2KXGyQIabpkt5yvlPWwBuOXzTu
uWpNOWclgyQdB2Ed/+RT/2K7MK1r665pPILY80HGOSwwhFKfGLmWJtMwd8qrb5mRMsZ+x/goLu//
zsFhW2WFigH/JRxkjckcRXd73TiFE8nVEQGuq7yr2GKrq+ET8nEHQtaODOlHgDqsPeowk05S72ah
TdRy+RJ2MUVH3Y0g+f/sT8y+7OqmeOV49JzwSyz7bGzHJy3GSsohmDc9Q/X7bl8+wglE6jyh2F8L
KQMLUgy4XcbP3PQt4I+Ip9mU315CqjjTerI6ZGrtB+rjgPGvYlif/DqaQY967UnHc/bvmsrluZau
81lXqm3x3Hcpk9qta4hOgweEPkKAFWM/n0SdxIN87aZ3DXJ4/d1Nl7DdFn3s2uU3uOufn52jbk/C
jB2rgcU/hwOZw3w9do3KBUkYMDJrodcaq45RavXUAqBbxNhjR7Hb5UTNwqxO715xcmIYOmbHQqNR
v5NmbNfCdPgLG6Eer+z1I9hyvfZ84q3uytf3OjA5bHYeuySFnufKpuOZvU2PNznnQtVS6+kZgAtu
+oNUeDnZ3NTbKeF1bQ+GnIc0lkB5KrihMlsOX9AuAxwl14Rwe0NydVaFrfTfI/llveJW6H0dNqUp
s+wEDWWuQr1vewnMVvR+pohrEoxdUdAb0JAXFSJ/nwxVJ9MSAyiVHAE8IY67yPJEQaVYqN8J1ig/
ZN2upel+giAOtciQfDyvLYMM0KAgWP6jQ9wJskD/7ZeaptGQbYIYQRKsTbzyVa9aWrZbYP3jGH56
QigT97EmWlBJhkK6iHU1IkPVbkc3d+ucAMxU7HZPy5+c9FsJ0lc0Bt6S2slZWu7EAXuXsEdI41J/
2Y09SBZIcQxvheGYR1G0L8XJv4YgcvDpDYZhwgm4VMPkePPHh6vv9Y1+pv2DsfkmIjZTdEH01wF7
oYvGhIKho0pAUi7rF85P7mRN51gAC2KpbVSmbjXhUHLjjkZBPgQO7o6vUfK8NgwyNOQEKLNAPi53
LXctnPRwd6d+3GZSxJTGtpOUU21ZDdkMUbKwd5vYLroNMz9RzditZoRspeyfgqTWAlG9WmYMAXwN
kL6Ak7LzmnZYTHwQFs9C7V5tEB5CVjnrEA8nWA8V4G85mQ7/ibsO3C4MknBG7D5CSAdAe0rPkc0L
l/iC65RqkUsxgsd9+PiSmeVoiPhb/bh3pYrD/nazW+aO/QrKiXBBP0olPxd0URu/3bJ+GY0LZIXv
VT55nk660MvFuIwMUfDKHgQoNklPTdWqKi2xEFxC9dLPqvgHwMUz1KBeMoTcSNpo1escpVF3ORuG
c0cK8hIU7TA+IoZpGX5UCjuq3AbsytcmE8rnizOc/jCBSMAOUcDaw+SAQIgIkE+d4bXxI+4NZC2W
K0uLuoCNa9hHs3eIC1A8Ollc3ly49DOPz8XQadHAbPdI5sVJTTr7BC80DcfzU6U8JJ2ZGZjY/fJn
obEdVkQRWxOX+VubQajCLnY3OzeNd3ipATvgfER63WTAUJg5WkmQ5NASiusPRX+O5gKaaHHaZOlK
Ivtb9cuPW4H7aqr5x9B/8FgkNBk1AJEYaKXicHnHOGxKLCyAyvCyunXoWGqIy8uRTrYZtT9c7RRx
mfnHTff6XFUzY8tR4xwtN/+Biz76XWys3WQOFijFNTr3kz+OYunwO2bnAuIV+w006cV9scK/NnSo
n+FO7+RqZN3hyugMsi7v1zzB8lJ0NuVVLArZJl1deAs4ko1IKURAbBNINgPIINJoXlRr49reJgd6
N3Ultg1ytS4BXPMQ42vxWAmOXBYKAhzZ4pTweSLzVOj/Ti/nFp8iXceEUooDzEnu8TZr1ibDwSqL
miKZB9oimfVGtqjNvDeHzZHJwfo4/tDspCrXICgaJKlUuhBdW/sA9J0qoNMnEpQ1C2B1IIeGRENj
ukWOm7zx603KmFHjXCghtqO5MMzK94E/qoGuWcPQyaPNVtwhYgaLcpDkzWOCRhwI3H1LODP/sLFD
1tyzSUjDpY16SoP4w15MurfMo9xUPkrCMi3LKYx8bZ+Xn7V5W7fL5VFTlXsZY9Je1kkbOst3aIFT
KRcRK2tFG+Xbgh64S04ERXVbtDw/eE5t1zaH5AVrIUH1f4tR2Fnvx/QgxAbvUcJ5dWYqBi9m218a
TuFRX4htLRR1aXzhsU8n9b3+R+VLDrYB6MMK+B+EHjK6DrKW1sawl6yDlNxm1gPlN4nbLiOXRBgX
sLGVyKMJs1Rh6pCwM9FQsJxUKdBkGpzI4XBrdSls3hPvF08YPFayw5l/OHhO41e6pB0bmky4oWqd
BlQRsc9Udolui8TWwR4j79Btw8b0DKGPUFi8vZEdRRCPvs9j1CWX33S3r7YD16c9Zm/8vxgx6UZ4
Jc8MrDRbw8wJGoQumki+jHWJ8N5XsqzUJq+2A9BaF5EE2XbwILqu7l/SQ/mRAnausuwvsNksRQ3I
aOFRxUmksIwPB/DJHn8n2qaFs9owTTc3Is5trH50aWSknlhfE2piEZHmPo8olibK9VGvQrHPHhq0
74sPZ+XUmtJ627Ng6TlfbMQw/z6zzWclpfjoWQLEyCki2gaaeuwBm+QY0jcpsFP+Perky0KEtApY
SafB1hQjbhGIpcHsJj2siuQ9RP6Gy1WxFEduv/g2cao1RBFAzn2ri9mWy/zSfcfTcUqdJAsqgOWB
E5/ClCXMfajzeWY5QQYqlC5ssMhL20mHwd7cb3q4u7iVOHBouq8RjI9UEFCGyOUfW6Mjz9bTrrM/
uTaJ1aw5t+xt4/msmMaK//EzZ6EZQMs/ZYQyos0+GIV1HWoHXXOLccB8rPRzLT8SQjDC73lsMiE5
8zLUOYY+XJCJbIYymLC3D+LFkgEA/uaqXcNeqGGd+zULEgj2H70z3V+qENEWJ4biIip2q67j95S+
/HIk0SyuA2aC6QkNb/Gx8tcTADT4A2IvsmXZqTtY1TDNZnlTjCWR9Qy2rr7yWeoh/Y1y/ES94ck9
275h6M6zNXeAsyR6TK81oS7BYOl6zs7PTzSYyP2WhlmJepYf9H/khf0A79h452PfVfl2d5NLSNcd
XNdJX+9recsZmdxGuYmsfun0sOehIb6QhxVxUQZjzWKossTdMevbgMhgvFwUgxoVT0KPA4iPcLyZ
cwrvmqJxXQBTPhHtuqzFvr2fOmB9EQJzk14n6Sr76m9RgGar2IflfmdU7RJQFjsHoDYhgSt1pWLj
4ucQGIZs8AnqnDEa+yTnuVn3ojRfmVXR41PrisJTrossaXqidycBnISuJfkc67xMQgml4OFLKH73
c667rXgxvkLLv93RLeEHdxf5DFFaqNWcKVMNpfykB9I1e2Ogjbo5DDTEa3ZDLY+VpUroZnhZrW1y
rpvMHwDH7YrhW8SUfUjYQ3VQDLI8m1eFBXF2qaKDcrybDl8gafDWiCJs1lEQi2Jjp0jrW728i8fy
DQCk8AJ3B+AfiZB5VAc47G0SI5OA7bXg0yDyii+Hf8SSNJXkkBMsqFW2rEvMA2t7Wtfn+LhXk+BM
fiyirt+BEUEUI1FkmYW0uC3/8f0gq09XA62HhnVPEO4XNtHnqJjr4BOXUK+Rbm6hLNGooohY3+jh
xrbMx/a3GRH/dK6BPX49J+kAVIVpqDC+nt2I6L3ojDQrz0MwwxD2aYtLe2bOus98edCLDC76Y+sO
PlhLbsJikxeTDXXVBaouDMa0qUdNuvSTkSVPNMFE5kXkF76b9bxSUeTR52f/gDlfTWayhlGHbHPd
0DEFIWztaPqRAytet/NuVi3rXD2bTA5inOyB8gNkK8ooEYvoQqTjdL9VTTBYDbUyA0y6owfWIZoA
hI8Rv3Fa/WzzcPGcNBReZedogVdiUZMaK4JqXyf9X3BmYY/lL/KjdkHE5bFUGGTDeUl/hcbrIhR7
QNj6Wbi9yyx5yn62XdI0twD7wbTX+37JAuCWncHChIvVTok5P9lVu7suxEfGxX5zjH90Bb6C6kqV
FtyGYRQpx1FElSpH4qZ3n8AwHWkVh/OcxxUjutBeuPzov/cQR38NYdOKHqdOkvtc12m510jPUlKH
WAlngGfgkFrB8nK+qtfWTkeroDR/bA7YT1+egV+2mBc4mfvxl8ViWZ82XLc7AErc+LiO6BTL/wYc
KyP8UjZnyhfgM2o1Qr+z5D+l1PKz6tuPth3FSPDKkH/mcvx7ZtdckXoHr0XzasRwNjqxHeX4deXc
ybe+rsuWrrDeiFTC7Fdazd5+NLHUZhjfJrlKTwWxlRcu6Kod4/Rn8XHGz5jy1VQ/b3V7Xahji5Hy
ej+NUO9cbNUjhiFTM+CchsgnFCMZuA/P4JUXPUFyptG/frYCqwknE1VE1XOprAW1GBVyf+heZiDN
uXrqfksiWZmsZ8cmju1BWXM85UyInMwZ9Kmb8lNTlokBLeptyYsHJigiFNyh1eLIHLSKflieHfK5
mNnEeBRSgU7oWPYPEzUd8vlinOeja5QxzJgP/dHGY7WaHxZbcuuiU5MUVYg5TDA/nonr8O/pbB/e
tDKNuQapQ73KH/IzjnYeVw0G2nMC7syO3RZf4XDkATjvg2Q8ugyIQXTNWS/gbZyZjXo6SoGXvr8I
vYBkfqZveziFGkB0nt8SVCBAz3gmTsB0cYTqMpsffjbLyAN8ucef116pJIA6J0O4jkgFDsXqf/EJ
WbwzJSUL9PxTI5zwZJHoWw4NVpsVuO5cA2AteSFcHvObcIPWA3mRtgm8RJItwn7X4i3vc5i0tZ9x
is/DE2ozovyJZ49gSnoiQkkXq+omerLLvZvh4jTXJe922i05QLOIfUBGwx1+lB1FY6iUetrVxWj6
qmPdA7dXzau+ktyxb9g1CY87zzlOd6C/rMOit+6JEzlGEjY7Iuk5JsEBeFkDNHJ12lL27sDsYJD8
eKQkPB3mooq2DOk2VpmispJV48+ClqwlLi4R4u1lg6PD0Tz8RVnFo9iYufx9WZvPe0uqouRlSnX6
Lj7566HqcR9m5Wl4dej2jtI8FDUEfqdGERE8F4GhP+zsli/xo0+huKoXqcwP8LL0f8B5MG1fBeAe
OIEhND3Em1eOEu+qy80q9AfutuzSzyfbFeQQLjErzUbYxFLqkaCmBraEPSTHzAV8BljGMuqLyw9G
Acbje0WkN8d2wQswmB6/AVWyc4DAFsEL+A8J6tRfpm6njwBSweyyUajDIyaZF8XHs3uN8a/1NMau
SgNWogyukAStG14xmZC/F0R7aW/CmQlcSadl/YNHs6HhKLhTpobfDeGXsTaHk71Uhq2PG3qltOp/
hS+Y2pPfzEWWiF++ZR35e9kh6aHbCjf36692MCqWkvwpscw/U3u0tMh1eBhWEyxOhWruSbS9BggG
1OugRUkGcsu9d/AqF7mSN2YOvilNfAbsl0zymA3J0fle4DNQIuvYH+FxV7EiorO/D4nnRQLyr6Xg
CtrDlFeqQEJWRKb5FXLh1TpCR4UP+CiRYrzCDNu/TyHm4YtxUlqa2B4s3iXR7tjQGojTFdyN8Rke
Cs6hGA/uaMahtpYFX4vwAnTOrl25v1gAH/4hJ/Q8uLyLEUpFZiFu+xH8ZtvH8sy86Sewovu+Urhy
lnQxb7I++fYoS9iovV5li7JLVLLupwH2/GVpnbbiMlqQveR+PsPhm2UBaZoPsZV+g54eKZVwlNCt
8tPbhbkZZuy5H95PfYHwR3ac7IddhxM6URsIS1D3wFu8bCs+18hwTKWoOV4dAowdoyXIO/+EhMF9
CXzUHPF/bB4uCk0K5aGNLaH//nPRRhRqiVWlyEE5uBhEx2sKjMHfq9lpimzqYpdAqlRc0cdgGuLp
N8uB9ud7366CY7sS/1X1/OAN3vy/YOu/STMokjJAnvr76ZniOE2maTLH7wMn/8i1qc+E9G3cdJ39
MBJm2MSlZSDPut/fZg98GGu4iokezXU8qes5ZyeoyIPd26eT7t54gFgIeZCTcytAf+y73GjxQomA
5OqrTe8Uw0Xt/rT346c5sOkmicYoHETrj0iJdiFqcEwXNbpkZgHRslus1sAiUamyo/06IZlCbmiO
/j1WfOJO+Nidn0//MXCcZzixCjkugWi2M6e1jOyVefCaNKoRynO6pp1NNjArLUvbtfXN9qYP3AYd
ezVcmVlZtgNH0kHXBjBlTId5gjIlxmsBeSTvKGudR7WjZKF125qDKMLVen1jL03C1HORl68FOrt6
Zciu4QPnZe3llTTd3q/L1BoEqAJbj7qzurhDEt4dRBi2c5UiRf4dyU6TWHtHhoNFniBt4jSICcvz
TdrN+iYw2+xGHY4BRf3s6XXMrd+8j9TvBtSVAihTDa45ZK46s/rTaBypfPPBeThBsXt1H+qoabVZ
KDHrhNFq9RVGXefNZJGVftkd2Ws1OBxYkZsd8howNv3WvLEivKCYYr/JsifWkJVvK2KqojQZ/IsX
omA9oBvNXDlucZwFlOYda1Au8yy+BP3t1hn7+0e7A+X3hil0FI1JzWdpZlMFa8pyei99hD27+rdf
Bm28nYtlKyAlsN54ipIC5uDCqOQaM3ocbiEpjnHbRnL0KgxvuQHuf0+WlC2JOYonHCZblqT1PhiU
m4W9FBSX7Vz45mKnkhk2zlrftq/iY0DJ/TW2g/dWG8S3MLHPjNaGvbQKIjiiKUU74eK6aNAtMMzq
tqO3LUs9KvLGiTIlLRRhw7CvtstBBw+BDWliUY7WIxnXmeiOh4f0zvbmYI2l6Lfx/rk+6ahWfo5Z
XIdvxM5OTxSQLr2p3zkzIoKbJXKTFqy99ujZRcQc5ukRafVh3w+JDaTz4LWmi8AlC7km029OfAYs
sdaenjrikAlWwhE56gO+IDeFFwt5TrAbQTP6XV6UVBiQvVJ19yN86R93O2p6Agm9d65PWNN8yCJs
Pq/za7TCCv7Yor18+bmS1VNkRlM7RDyXBQmvCO7DtE3kbwmAnkEb1MwSZbGNBjJttxC1bG3I1ncY
SeXbY1OwI889SV4otHo6Hm3rBpi+20bYZHG/hbODh3QCrj9gq1ajNfm2QgQhD6BgzLDJeJ7K2hdl
oEKkpe67tErXMY6HFmPFR73fuUkX5q/bNMcQbSpUOtLPD+etiX2tAgOm6H7mBRFGZa23miidP2hi
ToGQlG+2nHsogMQZahNzFCnprx8M1VtCi6C2w0W4trRXl/7uCJDcjcR6dHIPU/mnMldPVGpQlM2m
JHTOc+Cm1wGXSGI8rnBghmRQWc7hd9encRHnBTKIZ52VYfheUX8WW+2XeZzM4A+NWazjL5FaneoW
InteOPlLjapSDq+S/MrU3pr0tlQGhxEAvSO4sHH9FB2mDomi0IRXYnIraLbYV0nybSej5DtEqpaW
YGXSzp9T1SScG8VdsZ/3iHqm0coKu3HlkXqAPbVll2L0Ef71H9Cn3cfoVDJgU2LSqi1PupA86xwy
wk2SF934vMJ7nBQINci8tkni0/M/h+SryVGM0blasktT2swnnJdn5RMVrbuhmbCGBqXoJuGcQbRw
ZUbxwiMGRalclEne6Q5G/3l45sk26Bier2kEv2WHqrmxftPIUxm/mR4UQWOR04AhenzoJCoLhuRg
6NRsS8gn3zxgNZGGlUA6A0VkLAhep3OF14Slz4jJ/j834SaQBK23beLUPCjG5x027QqWf2EmVDwf
LkAan1X3pxreDDLtR1jthphsasbaDcG7y+KDvAC07Nndv/kI//ZI05HRemSoSDzCvKHjOGUdNcYv
lqxkAwK4CkhxaM4RuAerCXbww4sCjzGasL+BqsswfeqaR7iKLPvLm4vMgkc138LEo+tFVFXb3SPc
ojRsK64spwA+om/soe3hPkh9SMw2xQoulJe2mnvY8J8aw4wRAOvjPI22d1zpSyyBytSghhyZUtX/
Id5SprJLjXP/lJsH9nB7ChEK/MhUdqc7XP2E4Sz8qbqRAWTpAO1pkuClE4zJDHP9O+x2LpekWW/w
eY290FENAZQOzrud7TEhJAK99fU3FdUyjm0v8I+bncnjdpktG/FJ0+JxzQeT0wXRFxfGUKdhcZ6F
OTp9no9p2EwGt224QW0ddNmM8e8nIbyUFY7VUvbjb380bGzFO8I51nxyTkQQkeMs7nTf/qng5Sif
eYixwWzLiJscpqm4BobDpo90zTqhtN5zVQ/H1JqbZJ6iaTuSByGOM1v53InKohrlSHeSiRSsj79M
HjjSskUaEsguU7oXcSdoBW0Ll0HdfUjNVfdqX8KuFvi/NJ8E7xIH5DRH2dZQQYNUzJGSWCJK4kth
3g3uyH9YvRbGzf73V8rw6+47/sAh6XVU++0oY1v1cSufGhLjdTGMGi1RE7fHAlHy6j87SO62EDAQ
4WCzP94MtXS1pnAgaVkx+0DK3c3XZPcvtjl+UMrXIeIatzvZe4nYlDdgzo/CHkzcHZMR59G3+hwH
dNFSfy8cBllb8RYS28jrRXcbAcaOXEDk+gBtrC0PgehI1TZzZrWb3YnZuOEMTuofoBbnA3ZdZj5p
ElL11iOOVxW/bTbikZqjFA+0nDeR1spwdtKMqqtbitM06n1Avf9/5fEpDo3Gh6FdaTxadk+MbT3p
T5d3Mak9G/84n0cW5O1bNQhdNRA0EOaE5n8aYP+R7ughzylm7IOzRZkAb51IXJx2S9rsXdcgLupk
LuVsBbRXPn+Ky8SYOemax+bPAWf1nHnbnaIQrel22TffCWNMoAuKf5Rl0128pf0R+vFlVOVhqufu
i6qgZeVvFIChjedYMnIg35t7EFyqxSGb8jguuTKgWVJF4m2tr+ODmgyRUXpOc17YODaCrwqMUQSM
yfniyxSnKk2tU5E1WbtXxWm5XROZwhR58wpaaE1y5FtXzf4a6ShlX4ZfySqZS8cNn4QrkFABkcoq
ee010F93RQBYCOmsSqrUIcjybEsn97LLDCle8pPoTmOWC5E1YbE1eCR7IDMPTOsbbHktnvToURcD
EYeO2OLZ7k7nrZf7mTzv7o2dM6Rs3xqesedoSA8oMVS99CB4Quf0gZDJanseOwANMdkSJVbJbFbX
+57SG2k3jR8lWMzvLVMeR0rlpuVvEoNK1xMYi3C603DvHsAPzubimYs8FBFFDivoTGUw9qU9Ambo
sHdlDZJzdqI/GkXLSWwffnaqHoE6PdaqRmdpA3XgEDO5zaSOPwSAny0md0PwrnuV0iylfp/k8zcR
W6+9IQqZz3cTR9fuXv621GSpcjoIQbKAHpaz4Y9j3FplAlb5x7cf2soXhFmlobQ629s5utNXHw1C
1QtXAO5/T15j6UsCIF3+SXKGe0mWNKrf9p6qv3oqFCArKuFDCB3V4lbBEBPYMUgSjkJDTFlsMWHS
H42MsUddkdwt2OI83WuF5V8EaL0UfTzjWoyN13FZ+i0EubAdpYE42vSZObqJTQDivMXdNkVJY1Ya
gB3gshOb23dKXFtQEh0a+Qh01V1EQ7HxaTmJtUfE0MYHRkjs2MeERvYgdlzUVMbsj/uA/8DQLihl
fOGM3QLzXziGHDvuGMnMEUFDCwKWFN9Rq0Rpp+8vPpjpBWzho8kgNiPAe97OKsiutTg64ANTsMeJ
KC9hrlLJbkL+tPI9IVPeqPkq49bCKYV6pDzVPWb9nDnGD8416xIEaqnk8fX1IK4AS9Dyf/ROEezS
Ow2R/iWoj4hlnW3KizvOY5eJViwOGHIqSO3s2Xoav4hFKNWMfS9+2bG+OE/YxCd1VRv7ecUrJpF6
sKm9QwUV4PmgIxOfN9rhenLEcjPwx6MNCMts32/wpgG/eNzaQJHJuwMwP6UsOzOwc556NmKiM0kX
U4/yL/IjDRQjmx5O5cqqAmnVZ2yKb0ZFFnNzSFtodIQ/9gUPO3UWbpvhC4DgJjaEKZ7ZpmGIfFCl
yxoUyMJQ3NLfoIw0JOTI94iSavvxT8DAdPIMFEYZXIdQN5PUt+LOPw/N6ciXFFwBn+ebJVi2bVRh
h/b2k1pyuse4UZKeCag7ZzuEo0gSbQqVvTwmO9zJwVWGvFhFSey5xZU4iVOEr7DnAfiNP2g9PzC8
xQcAmmGkPahCG1+4dvNn08SK/hxz5yKQ0OuyK4YVFa9VcCDUepp93TPukx/zmgqV39KXbeTIHS23
shFzOkhhY4+mNC/FuHYD0P+2PNNE0YyibwD1ZKF01nW3eUmH7hfrpMDlnZpBHMWL7Ua5RAjr6o99
JWZRPmftdqfaa1Cz6SBIL3PqQaXkTzcH+ypirpYOoxogLH/tZN+s736InXkDT+AyqCjNRxqXTTVF
nstz35H52st2w43mUaXZzJ9o5a2Cj6jGG5gmgFP/OEERW8Y8LHCjAEIionQntwV30wJM6Bab3atA
pQuX2SZTe50iur7YN4PZfwTRylyB9nDHYTQHLd9BJ0RAfdb5ZojHVTgZarGhVkHcVDd0fT3OW6Yq
K8Ry4HzGVGBDeogH3pUVjd93Mezis8ev7TjKoV3wiKkXugFwNQyTaD5SApD/XZibFO2ZaJ4yBsCH
6NMrc6LZs443Y9zFtNsHi9osMBKtDuWByvGn7Xv7FTjZc8+EPx6z9mi79aXstTeRbXdBPQtQdkeC
1K0hs2iC58xaBtpzajO9uBABbLZ95+4XxSOSrhJ9ZnrmxAOXG1Cz6/vPFzdQCdV4gyWMG97lcTiP
OQakZ3SWREVlDIepDLSUXrLIuXD9b3Ha6/qsWdXpCfcFOgOiTvPjdwew3SaiC19g5YFcD7YcN8vN
405PSfIGIQmf62aIM+z/0GRl0zKA8G7InIiWsqtBawdIlsEQ2yTQMZacaoVSEzGUE2Vo25eK9VQe
gg7PysvpVnhddYj1fj/YZfB7TsqWotdUrxOTpnSXkXuzd4CnWY93eDhMwVDptDsMGLcuiywZkGhE
pIce3pFwBfQlUJoKbD44T+ODLTnPqs5du68BZr+ZnMDxFAcHnev4kVfrVqaOJzcf7i7ZYzQZmHGw
NTbPZPjoZJXUJ+rb7DpwNqb5mN2IBndeevJXQgg69mAIvKUeOSIlMtr0Kqa6XmOBgZ9KDBJpYWP1
mlYhznDtiGRXCvhYsIb5SYTeEP6I6b6x/mGHmbFiuaCfnemgq6AWaRqJe2433mT4JyIdnX4fZrkE
YvYOpftUlkXgy0ji6CeJMSOLJ/zSvIyuGqNvgKlXDRV5O/CcV9xfpWmFpIrGJu3Bvb35Tx9MQzPn
FQDk+tfcULcCWxrLMYB12xf5b5ZcS9mJg8eBhiMndLVQOb60IdW2IUZM1/qUrgDPL4O7kRanp77l
7UqXVdmw0Lg5ljI+rT3ACOoyYg55ntLlM+EdXD2Il5wHWVuCif86gA3KVfRFsJ1QhQsWXdrF4HHu
/9+Gsk/X5DHT6xS0uVxGa4MYRXkaOtnGz6fDk13znOQxEkdOOq2/ab551q5JAYl0r68vK6v01TV+
V7vRPvMisNh94z7v2DtCaaOAwghWKpQabMd5OSsdw4mz659d77EVviJ+uu3GzwX9vELG/OIrQRoI
/YqAmejx3NrgzRDLcorxpe69IUYJX+11XibJHM5QLMPEuAgEHvAfssJVU/QCdfXhf3TbaeP4Zn1u
yjam7ZrzKmjqeq0vCO5DnNdD1tfDZcZwnxz96mJsQFHWULstayhnsgxzmx7WCA65LBfOv5LYlzKf
yHJx5JGtqFQyPs84VioPsgiKkCTfCPTTLnPmrgwRPYYb2uuwnC+HRU8mpzIvjQutL+IwfoZtgsek
tjL/7goqpYTTT33zRqTnC3VW4abeFwzkl+orju0IrH0VhyFbyIh9MG2hqjQt9PB8U4sMJ6YuFUqX
OZyjJBSCsl7OPSQQDPA1ORnDpCI7nJuehHmuI7XjPId0UJv/KOwc5OC6/gFhisKvHK/kohvMUkV4
oIUeZvfgu4kjSJpvvK0iugIyX7GuPAvQbzrELO5AXZ2k/sJtAn9l+uw84kjzLbk4NOrDBcRieBCJ
Jtc2VyTDzzEJf70cUFur5aQ0Z2n4r0uC8ta6z/ysbpsk8sgl582gmDSa0FmE2/e6UrtYxUaymMpl
prWxZa5gZK7YgnNk7ZoN1ZR9g1iJxkSV4foAcO1oVayq1uJRobnyuJ75Q3ZiwBbEFc0hqkNcwwLk
2IlYp6hcaXNjZBd8Yduv1m1xr4tYFtXaJRT9pVsj0JCH6RuAUEn2VHPOgtAh+CufIRBZTpierkdn
RgjhngIE1Y7UYEBuyJ/kD9jkJDgtHRcpXbZl/wCNUdHLZuzqD89T/k5+zoDi0NMRjpR1lxpz3XXI
YjO9Dh+eTFqFxKcEZziyy/+UKfu02HwqcZhFNOHTvF7eRFKrx8tNbOTm98pnZ+hl45G+/+IGNaSR
NE7+oEuqtTcSv65bCUYKFByhXYfTy7jx5o1OgiO5AcKYYX92OQlOkgVTjLc/WV2fQFmfeCnjlIgX
I/HpI/30KlnaH+t+l1G0q47poP6a6dfWGUmeM4kPssrk3r6b8LDR56KyXdXwSUDqm4k9ZUTvcVZz
GJSOQBCqPpN41LjMfqA9VyXUkYBNAM8HwPMNdS+6NSLhqKrvZebn+Z3cJoPlp2ilwlIIt5/VoAme
gsSG89lpG5Jfapk6Nhzn9uxz88if5oXa1MAl8Ju4XMr0BZf5NaJXWlc6puf5/9YhYIHR1gMouCuE
6Kl6/adLCq+fh3nU9j2KopWy1l8TisV6iI75+DuzPMw+KYjjb1/zv0BIDoCYFKidT01ni4OkyXoq
NM1vloIWpgeQPYk/9VcYHK5vDI7jhgilwz3KibjrZd47lvIFzqoGW5SA0tIAfv0/2S2NQSIzbhHn
ZQaWtDo4jLhJI576Me7C1L0NxD1vNRhCng7ETv56pj5QapMZ7pcx7CDe7vGhWhkrtgTQpWjYi+uH
lrccmgAnHegGxvqcN9Mz2kNNXzL+eKNcaEeCoOjT6DplZCdstLiy/TSAHK2WIjTyRsdSdEHWN/Ve
+O4VmcpBKNiH1gFvBx6VtJIbpYpa41J82Vbso7mx6Fgh97HdsAZ8CmwsZzFVnab/Q0fnZIiw5QoF
QC26AWE9q8A6o0Cnsh3Lc7Iey3EI/5nuLzVLrg9Xy5v6AC+A0hWHoNeltDUeVktQkkFSZIPXT9CP
sfONbtr8EhraeuNN2p/Zo4PNB0hIxmUt67WtiQvaETMlGRHJ1LSplMJTFX9CfdToQQjeQZYNLSM6
U84SsucdXt/kTToi0ILU1q11PlLI4JT7nhqX22bxonKy7QZt+lRP3oLQLAmVkhflbXBlxDvF5Jcd
//uRAbM5x8/eZQ1VuAmpE+JijKDGJoV4ss5/9U9S4Q3uPsWahynfdaRUZfxFX7g/Oa01DXFfTvRM
Osbaqe8XQ4OmEMTvhWGPmiA+hKXU9bsFjiZWMK8US/5SbBYXuwv7yqha3+Huy3+wUliqMaZM+4Ll
WerhKQqJ9Se1BkRYoeoPyMmtQYQ2wkwaeWU+mzWvcYx5lGFTlv4tQprbeGBGIsjHGBa0g90FicUL
fP52no614+WJ1EAx+xV8s1rERq8clXW0Fhk0GPdrj3bBlJuiag2VoE3VgzXu2wR9CW3XdhhZhv5K
2FICbXAIvGIVd1xRY9JuHeSaeQJ9SvKNntr6Pexw+3qYzGxyLIKR8x+GR1WqvGvNQEUxdzYq/amC
a9wQf5++m4SAf/S8xzLIRrmBsFMt8sFXTtzqscX/4ceu+DhNQTDrVSGI4GRWAc7tQhgFV0v9mH+I
JLVTb4r3aEBslPxcKH9UIGX+/Ssh1OUR6GS8YQ8dtqr/FCSMGbW3EzVvZqSB4VIFWbCrC9lhxdji
RIDfl6O/5Wp5fqXaw3TnnYwQhohKc0dJVluc0fAuoYyz6rjmwDv7NiU5zh57uG2FZdrpThYTAsZU
dLdnCZOdhTA6eB2RJHneAReoleHrd6wwrnJSYLl0KvWZwv5OJ6pMCQCdMEgF2Nc2Dc7921oY9ILW
0p0aWCHHwOKjPkDRaLeTMErMaBCBE8S6gVjkwOo5/xSblNMVayJdplZAlblqfPvT5W/SnaUZIbdD
kQ13Xyh3aS94+XZuedMZJeQEOhIDYZAnJTr0Xj/coMPLWvby6q3rA8ShTO7DHQUNt+I77VkYeao3
MbUTTPhp6bvkRZKw5QV7kJMU0/FskMFcWeSPuT1qiY2lXor4TOx5P7QqcTYhFqc+gqCoGuUEV28R
LnG4C3DNi0nzYpAyd/LJ/Twzt8cSAU7uS9oww9KhUrH9/wiQqgDBqIFH0PzWrnXKvmc2nyYccwRp
JxskJir6vjbgsf5Af6wznjbwJMtQmec2zXBg501OABvyMbT0KzQMefSJbJvFmrX8V9PJaIXXIIx0
/TK+EhvFb+GDlphaDQK7IGHWD+I5snwI1nz7eoZe9SJhc76zaSpqnXp07hslqg8x30DdeUUd40lk
zh+ZLSQIkMYIXXf3g0TyoGccvOQAafQgKII3qQsk9LmmtDRyUCZXCWU62zke1+5M5LeSZOLwRI1v
tjNTZiqnHoir5P0nkBjZTEB0xjKrLo0ZmjJ6m3WsMdUX+N75mCvV03mieaWAvMtmk/EJ6oJGaM8I
zyWsXe82CUZGS/5Ynwrskgo9Umps0UVopmzEiqFBkhYNgVQmQ+FgDRD3uFMzoptb9fKxsPMV5rpR
ubm6jCR7nf6sGIDcchPtx18R+89lIfK5SSYfnyr3xvOp0U5IBoW0Bn9+dPLtRWxmH7ayCPTjaCGP
wuLrVAfCq+K+BljZHhuMxPXWmeqxtDnc4xUh7kjXDUXhSUI2dlDjhcCDoCewEsEd/2xgW0lx1Al4
5bewmj5AtrYOt/AGTDbHEt51QeFvLQuBkBa1M5aQIX88RHawg4Ygvu2rAdabw/MHKQV6voYapkkR
a51HEmXzz/mLtnse9HGwT+gSe9bLBYitFZdK3g+ernhFlSco6NTXi9YlGusF3iAmJ+w1FtZVq7LX
dNdz62wKLEe12L+iLisN0BmO9UFaQRBiS3lp/ls/A+DBD4ld29QtfNsKBNshO1PhCYOe5bZmqV5C
re6JJHsJihVXxFiQ2rE5NoFknV7LBHpyCHBddk+u3gaMn+lTbcTLTkqj0yeebngVwJaUBVx/HpkE
ihnDsOGGehz8LYd83nKD96q/p2P/lV/gFpSTqtSzvcJ2Wz4iOB4A+S6j/ka5qs8RmTF+5eSY1VQp
nXbPdQ0SBlfZjIZacadsWKC5KuY2N6OtHtyxMgQV60PSDqH4861diudiYaWhBlXlodIok7qsKuBt
AY9m/xZH51zfJ5XRJGDNLLYoHxD0gfTKYLhZ8qM0r16ajMKqiT2H4sLKJawoKNQ3E8lPKhHgPxTB
RDIHe49aZuwbgeV+tDdO7nvkCEF1bSibslwoascchozWwB9A8BIFPhMkDZfIMvHJGpkTwrDfTjce
OqDbxOOe8ZEB0rL4PSoO2SMa4mwpSbWlDMHz/Mi9NOg0TcKozehHUC3ysAuJ+IkNl1URgWppbydt
MgezoCOSlPeOvrj5acvuJJ2bwwViJeBBpEED4VwtodfhIRbuqgqsq1wmsVqQQu3fWeGFfSN5Gikn
ZDEVfBLD/JOGA+TbzvYFr5Mkt3kCxjqpar+9JtW45RTgYzapO4kk6mWFrwZzZSyUhd/9XLfJe+g+
HVo+CIn7RJ0TfvW+i4h0xtk3kioMKTPSO+S/m74yyx1Vy0wtGqRb03BFDFkV9lNdkusWPDTpaoAP
39uux76KmWMKB8XiDTb79RXahkpu/0kKhT2jz1NMYQ975vgfNM19G7uf9coGMbjDfk/XJ50wgSEk
gdzWodNDxKS+A784+1GUJCVMVMhm0092yur8g/eYjUDobTsQzrxyIVM32hungztYynVAIVgD4HZN
rQTV8WTCM+Zv0r8qzxI47MJ+7vtMRCr7MgGlTL1NmyMhsfqCJAGCXxokQNBdJeGJuyBJhfxk3wgJ
EQHrHvsbvxxE5BELSkMN0QmvUz1Y45ou6vQcJrnmbXtsiP3YoVjCMnFBlUO7gKvss0tTOj/Si3z1
IuazUwf0a9hYBKPbw95IdPQQNBW3Jnep/Yir37cBxhOkos6MZGTyqMiChD+5MkpqltvlliHkl+pG
WreTb0y3F21HwpI2d5CzGWflOPIzsjLewgRbgcyOQQazasxD6Fj/XWLWW6EIezn+YzbIpesdfJ84
q9rrwaJypVw8K2eptW3Dh+qrZHIZxJ3OrOCSml8tU5cvKje3zMGvr7BACevYwnbZfq+KKT1RAPjx
JRAHSzRLOpNxcbj3++EkXqle9e6pHodP0RhfwI+m4ysxjQqzTw0lm5Pzr7zHVnxDB+eF8Fdzke1H
bi4YlJOqNnZyeuWys7ThqMDnHskvphU/jlgSPkOXk2+HeIAvPlz44dNT3PAWewaGeCzqcDm7SRTH
n8l1t6Zg5GTlstCiazZtPzgd+r5Qazux/iAB8o4YsR8Gy9tBlYbbTuSp0K3l1jOuA6EKk6bdwmoq
yWOWzhL3vp5rBC1JzgbfrPR00x/hjrZVQbx67bjWYYzZqwDyTwgHe8pHsH7VTF8SrWNqwTQjgRxC
r5J3JtkvM+GlA3VZQoKI3t+obBMl8unPAPmy0AjWVT/YcQNzlilak4Ur1hDoXqmYzhC9iIl0VGUC
pC2YuNjEx8Mn9P/TlO3rVobDPMxYaEasJkb4v9+5LHrYRyAp0zYqNTsehBhwVCqj3VSQQ5bKHP4h
UEPqRqXEoxIn/GL6tvdhXgBMa7BbCxB8Bj9s5Uxx6losk+J58GJMjMF1vH6vDd61vx+T2ae5gOIB
htmIjv9yBEoAlUvkGhmFgnLEUG9L5IjGaytOyPRPfSFymiA8BwlFCl410t/1aL0OUDxIaWRm6kTn
6XGEE+a+fgNl5Y0SLyWVmHUk9mhfFIWr0ck5BvYCF+/g0ZKSL3ncrwJHymd63c484odJNM2wSdLX
YiUHEkU4hIUabnCg8FBj7Cf1c+YodzagosTdNT6IKD+UUt0lR6H9CcgcCV2uaTWPyQ9LX776osVt
3T7rLLwoiHz359Ubq2UTZ55B/Yv2PjbhPrIrErYgUL7kky6/BurgZ0Gzn1bd+ix8RqpSnlef0zm+
X7heUjnHPMAhKH55Qq2NwJYcAF4cWtzstLdNTqWkN0gFBBVdY2gfrRpQIr+ps7aKd5djwXuZYCep
v45/ROiEr8GCkrljXvwL5ZtsfCZUsDIa2NZp+2CEVRoJ8jXfngVn8agMCzP9MjqrEj80sDVnpOGr
LxHyKaVHblwPGZ6CMrz2etJmcvGYj2RPjuX4ngBD7N1iCVMhQtJXkBQhemKlYNNMGDUiWZC1PotH
xXj71hkPGELmAkOEhTm4632KuXiYXmJU8EDDuJ64g8atKJFmzMCCSXtXK7fkp4R6fDILqS0lpG/j
XtxAg/uOJUhI9vxhiSRHm7Z/NPsQl0ODIqBK0n+ZpK9795RwbGNG+++FRSZTDcmDczAT9uhsiw4W
SgJXtfoPfUilEYwsnCPQFSr9YXZmXnBcvmc5dzX4FQek0b2x4+Q2FzvgUyZnZy7Nx5x7Wo8JXbJ6
ia2fsX35pi4SQPp+24dzHHPgjugTTXcbRyNasAx6W9ajNgofoFyrJ9iZemS4nH/a7ztZH07H3SsW
YS7FDdZ6RLo7pNnZfxeEz7A4gRnKXRq+lPGaDTsb09/o4m4Pe1gqjpJhaag98GZgJVl/O5rg5I5c
9enhaJO8TKnkS077vR3yWfZWVlJjE5ub1gn7uFIcif3dMxjcn814oMudzboO7qeN3bnUb7yTGM3T
rj5fwTcP+clDalxonj0bASg5GFui6KhBOnp9BAZdoq0woHzQPVlUf2BiKm800cBR367XMLPiEZPh
+u8c5y/jvxFcWdkHeKrXIqmYJG3KqPAho4pCEe+gOytk3dQL8uphlKC0EptMiOvzsHoLCkIoV3ot
sDzyld1PYq0mioe9YKAqQap6ey897oLSaH4A3qSxP0f8VV8dU6m2fpQqEZag0kVvqZm26mfJfqbt
Z5kEJMOuiQzvEcnQvYaBXmIPQaFGJOmjr9QiZOPBDUMDJdoU6S1DHTXgekF3XCgu46q9yekhcmgI
EGtMfKYXuNknCR0vCP1MMfsf1HBvBlyMEq584sw8nmhWrLvC0tscZFKheyKW0AHyTMN3+tozDHqr
H76m6YTlt+CgJ1laYeMC2Z8mtZOf/WHA+PhY8DAVto4ATxCY+0ICiyxCq5BG1TmEX+akEqJDDO7A
ZSqPGnrMRz4QmpkoBwD10Yfc4Q2Oamw7Z6FA6RY6hTmLuAyinmiT6Jw2/k4juOkzUtM2uV+HAUzW
LiQ2/ATcDINPLbkkQoifeKN6UwIRBDpDgAGGgaeuzd4GXyl3U3ibH6mWLBDoihbuys6XH0Gp7/Ll
6OsEuZgmGUCeNs/wUviwYWPsySbOc8BWP0Awfsf3B49oeplFpaKtnFcRyN7/dMIgQp20f1sQIohk
aDHt0sDOUbpZEZz74vJYpQxaPi23YCjyVTF+zGW1I4ArQiJwk6VtICmf0KbgHSwP/0SfhRHrE/6G
FGmDw0IaxwCoIlvBdU3upyWEA5paoGGfKgxEkHgbAKsz1L6bRLUB98XA/mwOt/wuZvmJEXaQumJ+
2fE6HqA1WOLdtE5HeKTvxL+A1/Fg+ET/rRi5+AJHMYImXIzniyfV67ziHRDOcov+5qRPu6W1zzdX
pQ+FZngelxvGbWXtRqVpI9q+dHfDdO9PlMkyQwxh1PVFA/l38aVFQNjK5TG2L36D1rSpFOAXyFQO
UNeJavJb6Xi5+KTUU7A1dWgfynEhotdG2dQK8alN4YOVM5bsb0zwTYgiMuB6euwRElv8B1cgW+/E
xAhh1MLQQQq6YJk4QyRZN/LOfKAgyg8Vh+cnonttWtq6NSAHcfen7Eu0d4s42Z2XnoS8SYtSnchS
1tQznIQmWJ9g1/wocu5nnpVa0Se8sVhfg7Q5bNyf8X2S0xS3YMN0y51pnTtbtMHRlCZ0PI+vtQhn
iTIzqM0dj545+tjZHhbpjM3I7BO6BgTW97qJKHPVoS4s7eW+0VZ38xPGpF72R6IKmQiuYInEDAne
IeiXV/6f0xnnMWZ/2i7yvyTTb+iVa24FXyMJQZ1Pk4VEF6OW7Hz0D6rUuCY/QsEStdS70DwX1t2w
0Z9s66vnYVuuozLSASwOdi5iKtULr2lI5omBHFYQjUDNTLrlFsw1tPWNbUiHg2B0X7BSDn42oagv
1Al28S857anoQKpSpOOzHbmZCqKeXclNxlPJa8/VVu1jqPB+XXn2usI4xZOBD7RtspR+BdEuMV3g
RXKSsHX0uLXBepcmyaK6Sq+LDJEf2paKF78XnvoiNhbFZ69JmALhhX7COKtEc6o5GolUUrnJx1rY
5tZO0pfNM9+Ix4+Vtjm9hopKgm3mbJzSwFHIEhYw9pLnc2xlnYQ+oKiM+ws8E8NRlpXpmf/GEzs4
e6jS3oTza8hc5SapWrJjJPbee3Nnfoz01KBAYOQfWzDxx/s1/X2xbXhWDhPAUbQNkLvx2DdMG4aM
S5OS+yTzR7BGLvn4J2gvGvCXn72cnQgeUJhtTODgQo2ZdngZoRR2vsy8O0JMMPLjujtKbv8aN0lf
IAGPdrtnVeO+PSaWWEXeqySZd/6yQd4fUDpSga4zotXzy6pZBGaZRHc7AZNmJgQy+TkhrowcAskX
buRevRHKhfGV76/t1bqRYg59RR70ygnVunrKuVEHYqwO/xjUb9ShBpsBwhyPAcnXLrokSS22aP1M
uT3Q94A2fG6dIDZ6G00Qhifm79YWL/JFu4l5m9x7M13hJ7Q2JzSbaKmPmDYv7kQnvGXlK0Uip79t
TjDERjYI3Prh31sqKf7lQ5YxMs+vwTEjc0SeuN7vpNAILS0gZM/BahCyv0HKbHYuxrserBmzdgIp
xR4QMeZkgjy3qFVzj/X6rFhLC6XJQ6yjk37SdE732CeJ2RStScagTGP5YltewFMfUy067q/V5SpJ
nfgs6E1VwzoeyjYClKfqxgqxtY2RHWZNVoyyrHCOx9mBn32fIaHOC5J3jomsDJnKno+BWZik3bK2
OowNMHjHe7SWv0vwZIIf4RIc3qN4qLB5OFwAs3ZmTPBJBQW4W1HV+uRs3Zh3zFdCzqwFmLuv8a6y
haSU9x+6hyTK6x8+Np6CPfdueoWOhlU+RsDMhm82WwMWkfgO4WxQgNguccs0/ihn7Fh+fzqdYPFH
sU4Q2OfehTCd1mAqnNdZAQO/Rlym6bAY8RTOpF5tHeMYuPFczFhIutqEpLwS3Phk0YmuMbC1Mp2C
keGcPBU49bee3bQ91F8nnI6xnK+5htiy7fXQmGAqqlWv0Oq4O/cOs0GxQY6tXBVow1QXJv1CcVi+
MvPD2lJ8u7OsftK7CGQQiQuGgCXsuLl+GDAKs/9tDBfy5mPutjI0ibOQAFfwzK62460qXJ0IIt4M
xy30WIgGJV1jZ8n6oHs9SvvkmiNTlGxaTbqYkQ5UOlBJAGgBVkG7T43uIHKQLclas+hHc5ihu5R7
OeRWjZYzEhly9T2/LjeLICE08xvGcSGF9IyO9yXI2ldR+cRlcTp6SapwW2Ei/YiXmi8s5vovLqxE
iFIiAwuqaQcAI+7BGGXjLg4Y/+ZZSJUMEb8NLqIfdqM4/Pi18s7jmGPkI8I1HXKley8XOZGM9kaH
SYCXXYzJtdZtlx8Gz3pwCJK3M3v7GSGjV/dct6Pkjts/wZjQDwfrNiQBXnWcnngZWRYlL3ixSf5g
+p6qqj60tWOEh8ADbiXru3MMAuVHE4EwpkyvNLaeH/83YcJgbM9ljEv0kqM0+qfcVWF9C1SpZT0a
ckUXMtUOZ15+0E1QmdnzwSgDlkBUfCtnkLKSc3XHsNobz4O9wR8nJ8CY40V5og8tG4bc1dprRYAY
gUjqFDtPfy63dmX+A/BFbpDqrMPgePz9uRTLFazLdIotJm7KAXFWJbRmwmV/QtGvvBwurb4uNWpK
2L0UJ1u3GC7Pxf1BB+MQDpNquTxhgkstNwlbDH3H8tsqvw4QDUlaL0DCjmv3v4PFcMKfr3hXkhVH
c72IB/40hqj9KeHnpORQ92NfhynIueTbBCvq75yesh2JDyuDq8jba39rhQa+p0bktKeNkbDRk6Hl
45CdqcKwnXPMWK0PC2iBi64fpyplRGG5SPm+e8gIB6GW7Pl6F9G+FVus+qHSdBJxLnh1z8ufVo3+
X7jjjj2zH6KyR1pkstTB7uggPuwXiaT7F34T2A9L8KcHHHh8kdmftk5EKYhxm1yb06jZ6rA9mvLp
yJQTgk43VQZd3sofNNa1rcsyzPb6PqCgH+7fG0jgdH0g5jh0cwHQMvMJHzpcT0CEO9OwQvwJnvAT
Cav86oYbkcp9/etS0ewhSkBdeLoWDRZ1zLy7sk02s1rHX44GGMEYoRHf1W2xAH32WUmkXBXM6sAE
xnsrjWZPxBR7nWsJHwHMGJfubpjnMflg52Qirvi8njhg2DJNdp3EYASVX4fFn5oFPc2HqCrGMC48
ROwO6ljZm70cWjQrIKridHgKxG7jvob+0bUw+32wotOXbsmkqP5OS3rWHjXmwI6ADPdKhQNodY2b
nFkPqMeYzYRbswXe4Y08vwnhRshigfzcp6eI7LBia/TeRn8Evw7cvxRKRBAZ8Y+OIPDsxCO7U9ba
glCSWzq65NfNaU8Xlcjc/21JwERig8OllUa7aIoPbEFNyHI/nxEA/1XfHpZn9alisJYsI0E5juOf
QLX2iQ393+ee2px0ajrRho6lmEPZY6tykUS4Qv3LKRugS3THm5Pwa2YHLyG6jw1Y7WlXmDCsndZn
yyoVsj9fY7qGgfIeqOIyGL0XPpztH0fNPFpkAn83fPBAAfU9dh/u7qEbxFlscUnpm4D4i8gBtkWj
aB8/W5ApD5yRL9TGbYkXq4VD5CBQoZVP/OerCbsnzKkf+Sqm4+kcZyxQfdy6IcD2R5gs2OZMLRiY
8LZQ1WcXZEOxKIzM9Cz9ZTdmPgDsrQ48Wxhv9IRkL2qnRmQ5ORjog1OELz3uxQToj6rm/FIdbyyO
zWctDBcAe6SOsbjVF0x2Fa78Fh8VTUX9gVFeUuUX462VcDNJLgq3YB8WDhNoqXpenzHjgR1HrEvR
moJMAZZ9etsV+KYN/R/m5vL6ukIzZJs4QqU6YdPdk+xUjT9LtMjbG8p9TanJGKnJO8xgqnxK5HFG
xP+Uik1KD5nfNONHm99sGKHXLx4bHJ/TBFJ9iOAhgY/lX7AmPSonH6xvapi4airDRpClge6syMRc
3dAmC1N3s6f7HQLBKfX4eOx/I4iEvDF4EQrMpoAlWVARKdFeHAhnLqAsRBcDapcm8e6kiEhywvdR
VLFFI0suZcnWIC98ibqtiWZjDLMKJtgZcYDNcSjh0NTrZ+x8+dWhrLcOadJlfNJJWekT+yGV195j
Bd3Ys65Lh9agAVxAN006z5tJaRaznzstyOyLCJeT9Ey4kqyfq3QdzZkfFEu0yBnkzG9Yc6k7hp3I
odNLo1mmD/9zstHpBXVg1HRkuxyCpBKcOoWKTSwLiFodtxV0KYGFYX1jAC97pPKHTmgbRYk+Qu6P
OctL+zkJoXxrXyRmB4k6XIVyQ13TOdJYms20UsS4OsHb0kKmahKjf4RaKhO9AZaHfVEINC8bDDbJ
KerDrA4pbvRj1xkSaylN1YZIglDh7UBpcshGG2tdJwHkhY3mQvT5wMyDleI67sRRdzNuWRMiJrwj
JACfTkEx5tAQLQon94wKya9DPKW7taVVpYSGb7Is5+V+QYkNHRMtdki6DpDl2suQ1CLnJaSso+qL
LptIQDDOxHlAxrqv2h4gU2KsOgI9y61qLPH81bhdhJIwtzjsVpXPaIEhMceljWYfQJ+9XC+5Q6yN
zno2Rve0oAu5jZSKcQhdUyzVTDlvuj7K/P3DegLcAX4hVRqjTYNTiUc7psFjoKdxA4a6WOUyPG4G
6JFNTR0pYlhl4MBHpORN9At8x7Ak+jn0qc5WzmyoN1N40yI7nFkyJZnXBrV4BmQHmG9Vtt8xh5TF
fjbv72PfjvmNXPAyjBodBeliQAwruptLSq67d0nKnAIXpDYp7RU9wU8jtF92Axc/Kf4dbG9tTIZY
aCuYmn4+JuEKiOPKEPF1jIM7QtsWLiAFdQOzayflN/+jJn5VB4Pqj+DUiayu/6zzSrY6X8s5Dew6
h0skvCo7mLktZWN72rvYEaUkEsZTSVj/5GvxlHep8oGAx4IUpwGsV8suw9fYFpIIaN3vpk2JztSN
IbiRMfy27dccfgzepYOtQxqttygMufIqJNNuFqMlDFasVrSzPaRsA4cjUOKmfX+6NV61mRomSDSP
sa05pSB9p+8AQ9G65rzLqxSCXNWjWl98ht/N8iPWya4K9b+Dv0d6gSE5tmbPFu4f/8HdPHfPH2lf
PQYz6DQaxEiv4y+3TQz9MAZvpNB14xVZCNYFF3vyhk9qHo43eqlgz3TNDfB599zEDRj6qDV1s2Yg
b39WKP2QV/HlucitqbtPe02205HMOAQGdzLnYAvdacQIGyZfExhZEtUhZoAADGepiHHD8AD1Nyr9
Rli/+zWKl1lYcdM5lKowY3PHwxFztIQ3Ni38H4A0GudEIxDQcB7cHtnNXZbvx0XQdaF/Q2NT2z2l
L/V4qopU/arK2CmaHFUKzOaS51JJTgNn5OYkzZvs+lhpe9xHRLit7LJr4o+bZyPD7obsVcfH5Kuw
rmQ9QTKYpqBu9CfCAoD01bBFoaaqXG9GTJNO5pWja1igkH0FJRmZjHaZpGBnvyk1jEyREwGGu1Ah
+QQ5mQBSMxo7r0fcT1knfaWlCCjzwedY9+QoZeOGfxkRdr8BfSV+ZNKD6otJ8KXNgubLcMF+dseS
QIR2TNXS65+ApKk1pZSxzcUMI+04mJF3KeoSuFNK/pTr0UE5sqmyoI3ZxDEHsKWYlitJIxcV01jD
y+OolXPZduBWiQYDyp4Y3JJniMDk7K7bdEmGWejAQCPKfjGKmC+UNXmrCSPskEHJCqTCWtWui09/
5cDJitIY2kSOmcX7kmknvnbFz0pali/UH/BOU5iXxlC81DjHI4arUMLcFikOnM076pKRz5InYEv2
qo8w4U9rLQkpFDSecgyQfy83+sbr11RbbCQEXSBZ5ntD3GOGedVMZmef5O0F661yTFaujrmbhRmK
E406OeTPIl+CpOIVhz85EnRe1+ESM4NpQun5qANwQ3ymJ3o5t800qO26NzTGrbyf3aO7j7IAgqJb
M1un/VaoJYIBQNWPzOgVXu6VES+XkcZjrv+yluxcvNQyeilYsXRjyAkelkGcFxQXRr7La0SRzZfS
W1Xi1iBY4/wGYJBemvlZEGYMvLQ1js57gzZ2VQB5zottxzUrWm36C1ribixG3JC12FFagcYqBuKh
dMP/3xdYQK44GhlhQSTocp8xAUnJ4DT8ppGsqDKCHRIzOLEM19NCoW+i9ElPZFQktOIq5MAbF32I
QVUKldgebvF1Is5k319RX/BNV1wuw0teY8J0nNu2oFkXL8VvH6PIgifzg29JPFJkmI4BZxPOSISI
OOrfWuRMTDP3AlLFi2OPDqAn54YXJuA1Xsr7QualeeWMh2FqttiKvRXqfJDgllPUcIqlKRmGFpvH
KjhnhqYpd4yE8J2RrUcf+JcyoQjAOoSUZyUr7lBLZYaC6UI2D2BPIvTLEwFh33vKLk6FUOPhnyND
RbIMCRw5efbHi2863NOg3LsbVNxMiEIHrGEwVHnailh6Po/f2Uspst06J/aKURq/jn5vNKg+Yl9w
E2m+eoPIUQKasXu8BMMVfhsQRjeULdNjA9HxYslZbdDDnHi19glThTSVTNUc9qpiwzoIXQnZaiLZ
HM2anA2aSPWDePvJMx8OfU7x2n+Snwc8xMYP3XNCiZkeJEh8prG0B+0N2W6dDEvOoSAb2Vds1Ujg
sccJMpPn/hEoPus0VJxne2JGNUx6oBLHYMynjy11l4Se5/0CLafHSQcFeuirM0DuK4AEyZGXRhEu
JkWmw3si9Gc/v/9hcJZuZWbjVA+F9QsoCsAR8l0opJ0dpd89v90l0e+EoSf+kX0SRS+Bmu9QxTqN
Cprrup5t/4XHXgWLRSDGBnCJCyAxxreibx2KQscS7/SifoJlAzEVo3qggF47IFTD8iBZ+q/Yz4di
3OOcF6yI6S3T9yrDxJWJdgXcw2Ae2eY3dDmiVMp+1j1cnrhvBTtY89i/hCVW7cNlmg/MikelUt4a
Svxdwvn36zWEiMiq1JhwkmF/lI/iVT9XuUYAcRvEG0vMguZlu9UebYAZtHQsORfFRdowkjgw4bYm
GRXpe1KAC8dt3IMuBXFkub7FBmmgMVdVo3lVx8tOR01LDz+ciTOyw+U6gb1a3RJit3Efl7mE6NgW
UpUs5nZN7yMC4V98v7DfNLn4xMCR7mfwi3jZIdf0ROrqed1cSUiQRviZE1GLU41EVID0yzen2SN+
hjFHiE9xXOrxzLKXF2KSDa8rCvfFqSEwpVKNHhxhW44zgbwnVxD5+x5wanyg9mUqgMIYqeG+3RpW
bQQlbsPDfNKkcbTtzhHiykFKeNJXhM8+snRD6dA2wvh/4bszh/fzFGYVvfHwjCXG2UWSW4fYzJkT
667xEi5wFIR5znTK7JCEVaH2mjPC/88k7S2qDk10I4oA2ZlmsCrOvj4RjpNy8SkCd8j83ofiKb63
U0nujESHVLKlCpoS1LcZDXyjWW/ng5763t64XZ0vMPE1/HUFLYr2ZmsLZlDzvwL1j0qUAYnNrwJm
aF7ou7Svd8lax6LiXHFddfBFijQa/n75oxK/H+kbZkjWjqFrvbDMM9S9ElKVn+nODc+N/yckC3qD
ooF6Co3Cgx0dS1cxyrXSWfdLwuJFEUWErW2e9BI+hIc74vA3Werwqe8RtCXCs/b6QoxbSvrbDrHx
qkaPElqipFgMFZOiAzJi3yFael/DxE4/QyaLUz7jRab3XcRISlqB9RHDUu6pAxGE4B3wlivGnCtO
azgr+ttO4Fx80QRpMeRqzVoYzG5EloZt1zrZ6VVNAMu6bvQY45tnnfCBG3I0b7DEkCimpcnA4h4J
HMrpig9sm/Q1/IYdPHwdj0vTuL8/29yL4VE6QNK3gV6d2Zt4jy2qOQR4plUTd41pDtxyWLXMeiFI
7mDJgkf/dA7T69RbsrRW6VfKB+rjMrwhBfOfBpVroy+t5xX8QLcobCs1iGl1X6Mo8lML/AxPu44p
RQV8C1D1wm836O3ykR8t307wPrHz26oKoesGkcqgI6VzlFx/YRmgrd7QhaKNX582T/ah6+f5saRj
BBnf3TrF5t4GWc/3g1G5WVsn4kBBRuaoRrC54n7kgbiskxwaxVdZlG85ywd/qlcB9yE7oNOK7QgE
fBi4KoGATM0556zds+SJhScmqLVqz2c0HMyczAQkXyafmExpByjG+VMvpTXfKyLY4IkV0B3pNtWm
cJO9zQrfUxgxHDPqSO793iBpsR0mQhRHrUHRR6BrnSZ+ql97bIBTavUsnGWI2S2Ce+LzUDBAcwTB
j/iWoPauPIdUjb8fcGTuDpejQj9j7qUBAKrE8MQLM9VK08Da2Oiiwd8I+sfvJQX+ppaomwH9b8N0
1Dambm/nRNqyBTmCAXgzt6w3JrP3ekngZh4YodTcmpXXlcB22EPYdGYCB+q68M5gamnP+CvacT+x
bi+wKEoLV3a4HzgamK7A0SmPzyAetr3kvEHLpUx2cjrU/Ddo6aGixdZDU6SDC0nkJLlwog9bSo0T
icw1alAvJF1pwrPGEIOeyGEhEWQ/AWRe+adJJGM/CMM1kWtr1TLu0D4ZSdp+2lqnG7kFyaNeFUQc
GELuls27Kxv+HHM5AxHfjGSaWSYQeH1s2DWR5P7YHTgm8wS38NlmhplxwY+t6rvCek/OhAWF8ohx
IVaMnNpJ6zkHoHG8ZpUx5fUJLET+J9UMbJ3ytbH4TfWwuWBlxLHe43OSReyc55N3EzgbjtAcH+S9
mSD1iff4HKEZMvbqD83jmp1iDy27fSPb6T8IXzkL+iummKgM1GVrMvqZAiUw3voMyzq+ZvekEuHU
CJZEz6D95TFQU6y1KTLIHz2O7KFMoyiv87PrzeIa+KKoL8dHyYQUMY3as5c1V34FsNeAdDuZkXdh
gMVOLSZ3P29QlCuoN8urdAAMqyMU/cOBUZ+DrCh8VB0UWdlfvRl8VsZZqSimMpheGvN8ldj2SLFy
UjmR9vMXNp2gHZ0YTKuViQKcm3j27xVNanchW6H3sHl4l+uAZ0zcmTr4Yh2pZE0KKOkJpu8M0+wk
40KvO5P/GyOfaX0/1Meuxcd0+EZt2r6AqND8gVVZsnzmfsUMuFWy7By+KGdk2kpVE8hwuh7gKej6
f7oL/VxkbIQlh8ur5ZBnBQkavGv0DJGeCuhbUYnu+YAKaJme8rHXwh9+FMGFJtQD2rMpDkBYae3r
qB6V5jPoeDZIMYtsfxsttYYkHinfneATVIduu6f6IbNoPcfS7Ax13qLoWikJaJQA6EqvelkOcufj
15H+sC7IKV+2wccGl9vbIn334E6D0wExm7vM20aIuTdI4Wee/qJTo/yTHMnIf9xgM4f4hmwTCwAo
jNTizsV7Dz3NBX809AO/v6tgUjjTE5d2rFPfMfGK6+s3CxwjTaYhTO+zacWxFDwAuYoL+bCFxMCp
VZlwSCHr5FAKjyEJPScOzBHvrj7b8HeEmcbmas9pab50PKP1hbMGZPgo82d4jf//ucb3Tas2L8T7
dkcekbh829AQ9GI5w9xW3A314MfvTDxY0z5lrgnOPJDaLQDaOsEdrEw2J35FCo6IWfno/JkQHAwM
eIzqSW528bWflLssKEql9FiCKpa6ehMiG/MTqvyMEUW7mAgldpaG4pV0j1uNiJOnDhjUM7Kf8wOp
sI6avE2egwkyy3L4H0HlRvHEjVvSN72xpm2+IlShpCqMK3HAJbS5nVWY7egBLRGdERdxTy6v3VGw
+JjBHLMboq7krri3GxvzJlaU4aWPXnRjKN9uQniW1Q29dvtYyVXHKw45fTYPCD6evDn/AbVhXFNY
ECY/eLxVIRwxWBYwubUjqplXA9rek2LcMHZZkFTR8j6FAozNSIr98h1TFcctGHkbI33V+2Je8kp9
RXv6aHS657O07qZurEBCp/DH8E5ztATmOUCagUJeuExOxJUuCWJ8p64m/c2E627amMbjJSgger4O
J9gZtDNTbucM1fCSjnvW1AOEDFWy7JgE05TBgAWlPEdOQIvvLi4AuVJMTtax+lM6G1fOvro5hbaI
irGPj4iJbOGpjgbi+2JSPwk3jMmABgQNAlm3hfJTKZg49qNKzGRsi9GoRJbQjGWIdiL27Vp4bKQj
gGG8EgV45rwbTLwM3X3ZSuaemm9+Uh09nZQH0gsF7/Q0hVTyH8xu+Fbhj07j+mgkaxS5sk9etVw7
3BlJ+YtFEUvw8HGdmO7A+uL8vGvdlp28b1oSpd8P7ZlziTTr2LiFo4eB53LoveQClzv6psejO6oX
GRRM7rIwP1kdzh5zBz6EMlvTP60/3gXyowto3XZ22n4Ks2JNHtXEDzGvdc5xQNw9QScjYyrp3N2S
gHCPFzRw7/QL7Y4lwQ1GQwgZq9LYFp+6PXfFCxLqeL1N/eteUOuF7D3seFw5qP7obEJPV9rc7QNr
s8RtiJmPoPe6tnqy070LnGvQXJckcISTWMRR4j9EElvt6zzKIqcTlFBD56NcgwTO8/WGFPpHZkTZ
NYxYNyCN5sJPsRzKmghqZJAxy2mAZmibW74O+IlV8egytcxQdzpGvMzoQOSzD/CHKssT8yPzyvqw
pOxDdPnh6wso+855QgQdROsYCyTA/Zk0i7SkfaHbHKwcDeTxyLH3KG2qPt5+wUhGBCrf1W6kVQCb
F/SsGeNpM10U058e5te/T95yp9g85V+CxiQzVZDLOcYiwjdYrNyTlcKsNvsg6okkn+HmUZBcSjmq
1tGh82r2Q3uG815e/afI7jf5vw9/JgWO+HlxHUJpc8EC+miD0GOQX2sawx/a7iWVLdfLweh+6JF7
M9MOlLOUp6zyKhn9NfbyystTTqB6Ae6YWK2geaQBIhgXudtjYjtw9uNLa37UqvNRWdzUiOsBa+3L
N25jHrjB98DXTp55nkJuz7Pl9Rw3FLodZ+cQ718tg1pSF5NQIgpzDEGU5mwk/84qsJfwsHbW7dna
7BAZ2zmAEn6Z0EUcZzWhSoY0nTv32F3WEA+z/HeGA94TZOMfvi8yDt73wl7uR/RFnfjfce51wMzT
+pwAiR1VE0yna1G2HfHOEYS4eV7AXSgWe+FgHMTxVfzF4brNlGgWxoKp2Xwb0g2aTkrqfJcXeKhq
MinmGduQqadOjmH40IOG2AKwyoOyw0yofgelXNmSLV4lHnUfVGd/Fx9S5j3fEdd410tXKB2r35pL
T1F4D3WM2ld5E9StH4A3vFXWDBX4nuGl1/L3Ql6R4mQrSifm+5k7efAgKN9LfoMJY26qbUJCYcMn
M550CmfKM8fJrCF5BSkzQH6NfUbQ/ZSt32JzgA0EHTMun1tvoMGb0UCdH2nQF6GNEoqQx6A9GXFA
gg9z93u+V7p/ZTdCRMnoVh047digadYr4INVH0oDPBb7BZit27E+SrjfSMDo7Y5waMud/5tMbWTQ
cBAF71Qig5Q7kt+uF1Aa0xhldg11q2LCwNrbjdNHLMqcWzdT2MnvKw9zNX0zeux0TFN/U3uLyPpO
uejadKWeHK3Hs0VUA3r1nrkHIENIXLbHxZGyfzehQLzlzO9ex5/m7y7u5AdzHo/TNu7+TsfR9Is0
I9dehlxx+53OL2WzBLAkrRQkb/xPR45V0KUk5aj7qNbjf1s3d55qBgOGQpBj+0m1BcGJXttOfO7s
tzRGhOb8l+AQkil+Gv3hd1uvaT1Z5c3YzM8TIEBsW2L/e5jdx8nxmKiq1z4bCV7x0oTaon51v3Ry
ZADcclM1I/Rsec2P2Fu5nl75XadtYlDSkXpyDhS9RqE0yX9ncemzuwuPwwIwOL24tkLcSDhOFsyH
5jFbogd+2pkMwaCYgWeWqZhJS8nL9N26I1g0GRFpKxC/yqSbhL83U4GvlPMAU1tMor8AAUyLiedt
JpxDNuX8KrtgppLAD1OwbU9z8mAF/sokV9Jpz+Sl2uZ9y0C4JC76p/j4VcDj0MXWbF9dt5CsYvBb
ZltwpaN1oZKNKRyFPECACRt3R73sFqWW/ojxZsC5Zmf4j2/0H5KPBUA40zUeqw6mnE0yh7WHSRIy
4qZjF+PK4shkpKaYhSJA6xMYv8HwqsdyVn9vJ8vf7Or9WS4JrUevIba6DDQJG6/4jvpI/pmCBBGP
YLw/6HR8zXUibJeQ1wOVye7JiYbkzqqAWk/B6n4oQCu+4yIr0mM4nbSti6Gm2geGrtws3H1hYJFl
L6vmxUCOjlWd9BuZp72bvhJ9OALkx9Z4uDusSYIO2lxpOYssrK3YkmBAhGDqI39bsrndkLto4hcb
SlZqYDIWcQTEAMONuj+YtT6R5Yy3INlehQ+zFl6ahfFHP/1r3+S/7jkXSpRYQMM5JFLO6hE2ZtRR
d7sr1bXCbQli0cT4CPCXj0RwkAKiKLQ3JOBh7ILFVPzLQPLftiNmHyNpPdASy8PbbW4jV53UbCoc
eFgPcVPzpRDf5YrExX2ultDNNq1rapvN2HeOxZKUXv0u2Am9cIxofhudhWVp9EUIC6l7MhQDlMIq
JrDpZIeBPxul3tm/vAHSFsKFVy1brTUdOHyPMvrN6aa6fAYsIpjZExGqJPa3qQfOO/Uw9HGhoDCx
vpI1nGb07L73kS0rPg5MRRrY3oEnOoUY2lbWIh9/+37X1rC8dlKVn37CxO4DiZwt0bd6Izzb3r4n
2+oU9DFLqEFFQI/sOihynLbUnLeXtIrUhQYo2sj+HMDhrkUTHFkZIZQac1E0LaEYqNmfbQ5qM5tK
+FZpJVfpMR/aIXke4DD7a9kW3+gFtklG52BwJKUFh0Jko+lhvWR4kv9ooDQxEXFwoAftCVqLa84U
Papy5qUp9wCdphZQDy2jnvcPQxuUon+n4duybCddvMJnMfKrYZUOdivG+D+KyAKonoJHzNNvkDF1
+c5J6vfKkpluxXnbthtJ436QYVOWwx/3SSJuV/+lXgqXmMUPEV+fd1ehfriaq0O2H7unNXEeZ35k
Qfdzq0Qi6O/RRM0bXJyVXnGPwkWg3Urwnc+Lv3dwfLFp9qALCkbJckgo+EZOk1OP5frC1bcMKw8x
xez/66XwVzPxaw9v4Y17AZJaWfXeVxWZxQTjSM9EWVH3N5rP8XBllSlbxu1w9q7mEzximI2Yn/h2
BigS0lB+bgoeT63FjnbHALtV+Dj6qkQVj2Y77QRI/HceuC8QVaK4lSUYiAjcwJ47n8F4073cQd39
P0jX1hd1skYh12BoBDqmKIuj0ipePxlKLYggmZQPOfm9FyRH00inQ1kFZuJnWIN3W2CubH4WX+IZ
qwA/2FhCWOno5cG9Bja7CbzS5C73q/qcQiSK75JLWp3lwEMPwO9aYrEguJ+aEADO0hpVlS7F2ySY
X6ZHZ55ap9AL9fjbi7vVnyPYOp4X0SkV4tos5mnoZxO6hTq8qnSHqnQ+y/Uyi0UhWfnvAzJPProC
u99waZ0OYr97uHIreHD2hEYK+XVbVTY1fwHdifafOwDE5PB9o6otgJcaw3iYqALsXSQ36401mVOC
zyvBIH7sh/9oZiN+sMOI8nPSSlCeqZ6beFjAUj24Uan6kSSFkEptRSFlq1JJ+g+d7QVDyU6l+e01
eoaBnT0bdggVh5wkPvTHizr6hFcJX2Na70BrX37tBjHIfEFwvQQBeY27QdaUPK1b6FXjCi5/T27l
gcnXQB4xLbkTzlLCwLpy9UXdtlcBXtyrO9Xg4jVg9wq46NdUnlWT+tfC4WngXcJgCA4OSc1sS0b0
dRddcbRj9qRjHNMYPvwOusOjxlwbILZnWqdYJ/XtgJL9ovIjNmJcumPhbg6T5ja6zEzOdcSTCebA
a76gCdjRmBGVB1+B8EUr+d8EVxx8/RFCu8blvDCtu9q39QgFv+LEbEzckfRRnubdy9JhXOLYC6Ng
+QoNd5XOh32K/AUMcP7ViilnFe0GH594qAFeloTfKvJoIwNP8xU6Lg6wf1kUrvZBAiH7c6CwDSiE
t5KlRJbx9SnA4ce3IB+SMPbxUPt024ntSPWuUyyYO2kWbRlAYUhV1MmVRnxL/sK1fZ08YRo0zhSh
S0uxhT8DRA3kxfzRzatzjAWlU3Xp4tl+Zx2bTngVb56Ju7L5MC3xJQttct9AVRm9Q/wVAHkD9rrn
vLxsNv1D2jeGtB0Y17ZBmVPmIms7OY7dDlAKxskpabB9saPFBz/N2afJoXvzCePRghFGC5GGX10f
2N6cPkpporLDSDfaGJcgLW/GkcZAzZ1Nbirr0aj+IaqtGFl3biFwVgtOQ83Qh6KDo3kAm37ke6N9
PspJhhUr75Af8OUEC3YI5Uupn9GInj1UjLJl+q9fSPiZSsZOJ/ut1OuCSUNZO/tb+dk1aR+SL93M
5ozD2rXrwQjhwiXbGHGIHwUgOErm1kfxdXZMAT8VgEjTHYdLupDI1/od2v2nIMAtBXHAOo8rmxOA
mHBu/ZUfjJr9OG3zTW1rLBWf7w00P6y7oiQIEAxZiippch+DqB87OdPT+00oSqiR67hUdNyEBpUg
uVcTA32j5XwBmJs3S+qzc6srlKq0uP1MZyiDkvAbLPUlbtDMAsDLszARgfZuMQ3OWTNISfrvQ9Hv
bYK4LhYclI+YrE+HGDkGK4SrGd5wuHRj6eJ0GgRnki+fuOnEzk7t0If/kE/hUO6HqVuvGaKfLdKP
rEdWLtpNYanpoGJpr2TFmMCJp7yxH/Ellxn0B7AqOe2XdpenYbeOx9rBH1aCEQTIO3ozb4ZZAPjf
UEG5iAYbwBpwgitISe35wF0we1CvsTda0WTVsLbzOuYRX/UDEPlZ07N4e968tuhnkvZWWvzV9id3
l7OEwt8xU4ZWreVmAIU3OcPnYhaZVEHHPVnkjI0gn2QXhBUeWYp65Vr83cikb9vSsz5C+KR9V3VA
OoqGaEHiAxK+k4lkcrHL0Bh5wX6bK5Rq0qw0rAVsC0JT61wGOFVsYYG4YMQTX4FVxkwUzuIjKqWi
OpVmy9Uk3hvAuymL3mV0OzHCUsFWK4MU8n1z7TfzFafLof+KQ2nuIFa8iFMZtUc6NorT1Fh9GE//
4JY4caAAymg55afILfkDx7JIYRTjcMG9NW/uOHk2xEmcRsRWdnOvoUy2PfHz+6/T2xbSy9O6+mzc
BkWHsN9qVJ+QHTwl9sNmJChu1EVYroidy0tWkzfvLKnqlLo5qPzCjO/613jCuDIolgqXC9TbDKkc
QleEJRB9zmt+kOykSOTeYbUjMPvz2RPPaxr/j4dwcUhV6r2y2Zv6fxN4AEj3EBrpOFmCqJVdlUxC
mWnACAwco45WEDiWcvCK052/14PJVthGJXFu6ttFow2PwwevOjsFT/C5//vx69qYV2iwez8HdvZu
QiSNpu61iqMgVGxouK5UXIcUBCploxTs4m2M9kC5B7VW/ULh0QjNmhU+duhvFzp6qbJI11FZLETh
xNhPrO6AEJ33nRB3HXWXbmVqk4x7FYmwTtXac4M/ghreeYjKXNAeuUU/f3k6W3RwmMrAiv4SagHD
0x2eqe6cf8KSo2M31neViMFlpVGf290Ea5JHquns1hf2HEVnptHYZcV6n32XOpF0EFW8ypGZL+2C
d11gD4m6wm2wojorjLoFnKp4qGlC/yjkdlsxSSfYTbv7ypIlw3sEZ89XhZV9eLo52CQFIpkISKVE
W3wE4wKynkE1OjuE4C2kNSihTGCa2mpGb/FULywAWxKhu0fP/eEpp3t4Z1d+Nu7ZWvS9gqfHDYZv
WIjvCfTdHloz+r+dA0pJkMfboysJGq2btuvLMQvy+qWQdV43c80oRecnTs9aP9pvGMJAt+z5ju0D
mOzhpcanxzHI7817rAePC7Cih4foapyCWT3cegPyVYf5GL3gjd5KwDKTrj092l/oPkBzSNpbr1Bp
uqcWHFRrC27it5Oa7jP1Mzejt7HaJOeDi+X9JYGOD04PIFsruyeXkpUPtN7dGE5hbUSKkh/BgId9
7yi+w1tFbgeqrtRrVpWVjUPhOhylN6oFDCXfzZKJ5icqpNPlh/JB4UfWPmYWdxWEYhdn5QClq+k+
oFc3t3zEvq2HLpP7ZrFemMMl157ckRZv+zOyDlozPAH5MYJiw2mBzyA8kGTZdOgkvpMSOFL9d+Cz
PIrZIGjb+obzGWWCcMel1ejpN2zS3a+cKfWHOnUHHksvG2dpgbZjf8Qec2awLV9ZUq9NdqMdifWe
MA84w6eveTQf5mXbl751nKNF6/5T3+h5FJHX723sG/IxiCkGgNi9wQpgBauz+x9MMWw1UWeucSkC
HEGshSord2GMF3CC9DArkSjjEAmsCakwkHtvrCQMhwefufFkLrWijiPDYRFsbHZl4wXB0YENvjPK
VqR85kHg06yR3Co4nrOI/hrneC7WyfD5vmG9Ew4cpKJ0GFuNIRc20x+XLtHn21LyRRC6O080QtKn
3fr6KhLpO0XsWqifPywedENFOn2rOHohMx36VB9xxNyY9EBNxRSOTf8WxJb7fT4rD/w+YsBHZ+DC
FpLydrQNnCtHsZhs5hyRlf1ufmaqQksQkB3SZr76XnOyQRIvBcloOICHTkmaAMEkMgQNzcMl6ScQ
yGi8/CFBTr6ecLWBvk1BChxNfVE4AE/04VppdXCaTi4XVs9NKJm6qXB7Zds4ZlPpRdSSRsXSwMk3
ilxTv1/4BIYG2Eho12Fbrig4vlnsN7prBwqLhghJZvb+wYDtezylp5rdXEoBOSaXDh+1O3XAr8nV
N08awgPgv/H13iy19R16QpxXJYqNvtNqC/zYwmc0NOFA/9jR3OWhITztNQkDcPupnb7ADuytCbBN
t5wFfcGM/MjAdVAvhW8TW7Q8erwXPWGtMxvcZbWXboTRq7X00sEsFuUqDSRVWd2ZuMXDez9KEhFJ
II59q5yCLSTk2Z60m4gO4xMaUdfEsGM2OVwg//FI0P2vgq897xgyb4qHQn1g8p2AorZjlCvsS56d
2wMUem7A2Jah6ZZtX4cK34oa0kGWUcFYPjs7zN/E1Fv/OSNTNWWdSzb2+31ymhowz0QK+htXty/C
DRCzKv1aTmq/J1MGKsSZUzoEgyc7/DHGPQOtsS2xLN0WwNDSF8rhvBuoTk4uCS7LmNmLs4HRoZJ9
7DpSnuOs7tKyxVW6SMZC1mxPt1Ei8Oxi5sCT8ZkEpWFHEz3oISBQ41G5trRJwdb6fNpf0YTbjUr0
ytEhRUKm06/IimjJTnukayPru16S4NhlLzc1eZ0BR914G7Il8rhi87Om1Dxc7HERpwZPUbJ6GBeb
iFdsg6wyzUefWWNr56w/WGQ40R/dnxZ8x0u4ms21ZiH1MTcU08mVbfph3mbP+8uGVacoA6m2Hnuk
hjxPL/XUXjkN8AfAnFY+nOMFTSd+vLE+XBE/ZNtM3SnV1ocQP7pJ9jNj1iSQHde2TzVQfEJD7Cth
+H17UnRV8aa/uimuKeKIG7qz0/O6fDvfxYSzU3y1Gk2r/1UhtSMnKssIdyvZX44Z8XpMnVSKOYNN
vgk918pBPh529CKaORJVbdPYK22331lCct8lWNki029X/H3xUZdLRXTYt1OUmqWRoNB2Mtxa3yzM
cXsk49Z6HI3dkHyyukdmKmlTJjZ54vXw9LZjvVxG7TCG1cuwF2o3sisgARSEGchBkrewPNd1EsXg
H0HzvgALdD986teABFLrVPNpKUexsJmMJkIyTdXpnGdj/tJiVvicRagY3EMDyW7s6fm4DN5BXLnB
obTEFCRgu0CAiWO+C+xVt8jmScMiHavh2Bno2uMFrd88EE7NH7fgEXjfnamlMzBRjsslN7AJMQgE
n8S8vUUbi+3vMt2EdqsPSYGrffEaTmRRaJTb31AYIyDJd83cYeFGq0HFkFZBU1X6+A0cu5juewXO
2Ec1qaUBsrrbYpIWeAMxspZ16UIXxyNwUZefltwfG5O8ZksDqqoqMc23u3r0Zmo09IeBqfKhOq2Q
dTIAteuiBjVEtnBWvcYebCdzcXiwQFdVVpN9bno9fkDDcm9r5a4rZPKbUza+EbRrtSASbcXodLxq
nivZFqSpBJZNjUFr6ZgatWDpv0S6nzrEVsp2wDPaczHgOEmqVzYDoEt334KebXiPY7MrGBwXK/Wn
n7ZtwSsxpxcO+9rCv1qYsGkOblm/FWHDBDUO+iI3abVw6VkLnqciD+7sFQHn1n0r3YzPcXRhZorQ
4KdBdAuE4Avb62sd/4eAshkLxy4WA4+5XqGmMeDzPRsH9x7yQsccJY0rW0THSaWw83duWOplhezu
usIDN3aAwhWkcmo7CEKANAssxQ0YbgEYkNwVK6V2aobqDU7m1aK9Epq7hjuSdv2JxuI3+IoA2PyJ
zO/rtfY7FZtb4xnctW5Kgu6rIk14q4Y6tRSiKn9zS377xzVYamAoA8d8aNVt/Rr0f0hAByDRXU4v
9ujF0jScMcbJuwKkOaIzg6epkTclD7kkvPd+6OGj/86HeKJBxP7n2E+IWoxgvZhNy5S+AXgYy19a
T2Sx4YOIJr11WvKzD6miYagkWsuVvZl/z6Zfw8H6ibw6eJhXOxE2e+QPeXeFAFVRvRReiDmdcueP
Sx2PWtQ9zSm+7N1qacHdx8tc8wE0bOSIOzENJQDvEvJm/Z37/oNf6tpZiL6tF6qLVSVD5FRUXf1e
n4WNnb6tpJJjVH1SUm6B+iniwM1T4b/9+oh2M06Up+NItgcHAZ5v6G4pOoNuylwdfmERVZ8zU5UY
AHshVgqYcdHJSMbLgJRMdFxv91l307xxnF2CPY07a0Lj9KDbaRvg5+gEoVbzyibBjrb0NZT4Fq0/
bwxUbIwhvfti+POLB+TVPD6wQK3+QYyopmi4Ipl4VqPNDQ84HzLMNRRXG/HEOW/9K+t8dfswwWDE
ybW4VcfWGp3q5E6qN1YYxjSpPivAYCZfDRfGdAzI15C9fBrwCTUuN8KDlVDc9Vzu5Ea86GCWY3hq
IHsnCptATHiTQDVdTArMJz+F8VNad0qnjlgoGOhubHL26y233qw73AyvmJv+9bb7Q+qu+V/iOXR8
QVoVCpogmVNy03nk2q/nvTf0bNKY6jHuj8erkZHOawhH76efuIN36ZEXdu3i/mEnEb2WDsMmVEo1
Wn9JDsdLYr2BgLvCLNUrLlczp7WhD1ydX35+inwfJU6vABXfGhV1wG0kX9RaSccNGqJOrm+p8Gdk
I6+THiWZBwTEyp5fcgJcByZcdTR2xNEQ37RcpH+mvq8YfpF9ebzahvoZMKhvrg4hZzHMMKJ1iaBi
JvT8acSD3Yixa5ikgNA/ynsfpu/CyA3cFJcBnr4db5gCqU5z7yv2qifTe6lvODTMJaCsF0C6UYSs
ywjoU7siAO6nBxlEMSq2CJHw3CGNIQ0GnnpqwfwS/pjXGhzLmNtNsff4iOBzDoaB2WMiW3VXziWR
tFs8n35nkAJYFg6Li46ktXo4jlv4qKZAY+6DSqS4qmxhfWMddFXr/fFkVzD07gUHmWQsa78y5TgO
+h7a5iF9tCFm2qit05xZ5zf78z10gJ5isiiKB4kboDB+gWCaaINuI2+68/9//HTica0IC0MXTvkC
m+1k4QaN6TzPlF0i35q9JIVqK1h7ZIZLiLXxYEIcOC621JmutjWVYgqxYr+uBb+MnNRMOYoj4Drq
rGno11JlviGVxaR4+8EdcagaGRv9nOMPayev0xNvdKnGa06Uz9XUm+iLFXnahdZHekTk8X0pS+ot
OP90apbTXWoUt/4ldmV9TvNkTH87kF8nhBYwMzSWXDcO9eoUjD0EQ6d34S0a2cQsgbNfGjwZzb6R
VqowzneVLzGVf1vLNqA6HYRZIp8MUOn+NwiMHSVzOmXKMpIY4NUPLJAOjKXKahcmYSx6GhxzRcOZ
rxUOxbxVDelib18w5hJjljcRYWOQ+Xe2Es/NK4DalRe8DKTETtv5BsjnSl6rHYu+qqTTv+PH2rHH
F99yoOnwAgQC0BWz9lh96qXDDeyfsdvPRNwxSB1yhu1rpRkpc9GgeVtyRgTDtEX8skS+rbqOIvEB
uShUOJwNnMG9ZBnEDpdVJbCBntAkOWOpnMVLJtCZAKngs3FJT7YJcmNslPt/AFwDVZe3MZ924yaG
u3Bx7PcE0J6dXDPxo5aURYYm7BwmsNU3q5Aqr97l35n0QeJkIsu1ti7lTXxvZnGGhCqQ1I3GxnTM
X8gu1ef/qGREzw4SoyR6Qom0UZmwYj56YNbHneEDczRy1ESW7br8f2m7X9Y903woBr0t8lVXDjZk
qNVwo/wAuFeg+Zd8YFnSBpqOKq4RstXUGNyJxyHrQAmdal4Fa57pbL3KmCfiTzGNbmxwqa9Ju58e
IPcfjs+cYfIcjpfVil/pPBGuZH1yFg30gfQL/Loq582XpEHBZdnbA5JqGbqySHuD7bYGJ4N0ZHBA
4hWvRjYIvP5rS/5tM585IwBx/ty04aq1EydGf/W2CDATxZR3la771FQSYTbmkP509qGNUXQvWOpS
sNw5dmeYr4oS7+Ck01d67GjcvwrbhMfMeXv8kEguY3ArHpR6MajmEDO+4w71uGYAgIvvUoWoBaS2
3ISuaB59pze8qjBRyl9VVM7aWWS+vaamuQR0K6Db0R3uQHsri6fft2yykRe/PHaGUpaWPtiOLYKm
mV7fUoZBEmPpxpGXmF8++5CR/nhqDf/aOoKpwLfxJszfDy673zJ+R8oAKUiP0E93YEKZ8eqj5Rbl
15MGZzy0qU4pOWQs1+89QiyzGvKctLOWNiPdJGReUA7/Lp8iZIx2Vuq1PLHz4NHL3FlMOWCX02Z6
gS1nPSgdLq6ieuWuk3KnweN/MqAqcrOp+aPFF8eCBMlUA9gzEWswV+T4Z0xv6Ume94gfiwA3Pgfv
fTCXcxPsSmrd6wy7kgqVszISgMFuNj0o1uNoBITCmLESgxqx2U/ZS63gU2crExMDWNU0/AQRL8hs
s8r+7kaPxGmU2dLZo8QWPPWegB8GCsm17lWy1EVaa5hLgvOAS+jvbyf8Q3C0WeYMzysRdpvFlSZu
r+YEkg8T83Rpnb+Tx6EujiiRMB0xunPVMQY5I/Zvvzgf+s9HMPKdxFl2WMYhzVQYILbaaTleZIXB
Sb8CMZM65FTq4ukrYOUgqptBZVjTIBdM92Qa4kM/XdDnHqBgrfMPzO0fBTwmexZ8yrX5cNtbx1OT
+m5vXLZCpzfApYCpywb8esBW3XO1teIS4hI2OnefRNxMcX99S0E+IkNON/nGvvewp7f/bMAWZOZj
H7ldXiv4L377ByAMl9rIpQg1hU0i/zaXsjphIURjqlRonrYTezs3S8CVdmVHrtmJi5KaoE8IWz4Y
3XUWTwT2pduLOzbv1ZPCfb/XNCF8GMpLGPnjXMRf2/ERswLkxZ5mRmu1IotVFyKvuB6Egy+vQODO
nsNpNSAIwy6ZBtatQHsqUI6zecnWoii/W3TmGtdJtBihpWBXE1KVRCGSbq22xorVGd6OQJ6jPu9w
d8S5UFydZKS7NP1wsRc57WdHx50qIueDMndSEitACUwqNpKQYhKMs6lGTD/9Fw2omK8PtJYQvUYb
RCChfgc+QYXfPNusAa6H+3nigvFd4xakNdu6p1Sea0BpXKfWa1tumb+swKI9wfeUMRY3/ghaYfMV
KNauKM4EuLmJ0Ps+tvtv61JyIMPTgnihP8CMXrBcTXxXNvM3b8PtLGBKy8rboCOtPoWElQgUdS56
6cbN+xbAgEjjWFrU3jCJMBvNdXNLyTdYFzpyH8QZVHMA3GXcbhK1sRnmG9EKAuMi3sEFY/mAXT2g
YS+VIm/7Gc8nbmien/PgPgSUJp7pakVrxJdyj604miEsvQ7JicPWJ+avJm6HydCtIUs3fxCdJVB+
uLoDAkuk8SwhXSVZVPLRhVTTjJdJ8uDUxZwugyEB85ser7hMeL9ZjEl+30euMTOoh4zRsopW8ZdO
8aBaq7mEUEDrDktzAHk+qy07w5YV7CaKeQ8+JJvdIq3VW4Bb8E3ydsppcR81gkjtj8QSwk5TgHsB
ZR8YukJcB8IH0OHzwRPGXoENPv9NsEAFeV491cD13LQ/WX+6oItkxdlHHMJJw68HAu3AQ4h4WDOY
cizWuxg4dcawqgfyKKx98FYzsfgOcotE0vnuxpCcjU0spC/mEAI3d9C4IOMMCW6YgCAHgnLzuzC9
M2+EGqT1ngDlb1Gdb6RG7/3XeumHo66DLSpID551OEa6W5v9/Oe3An41QJMopNmDfYZhKRWOMzSW
sfweaRFn/SY0mKDx+Y2CYHLNCXwOtWFSB917G2+c9xAxIu7JK8T1SPieXx/m05WnGhwC467qlctc
SySmKCer7nTUEmZT3Nu8QWFDv37t1Lpk3xmFJFXSrvEUgTO4TYH6JbbcTAWJl9hqtCUcUgDamtvU
SOd/x7rSpgxKpQWEB3nCTd8x2+Bzef0hE5ifFDvLQNK2Cf5jzPaKuAdFwJZXkFOsk6lzl0WrMBgm
C5oPQXX4iGn3maaCt/nbTxt5oWDJz9B9wtDbBJJMfafWe9HtQFfpbc3280Csule+dDfjefO57FZ+
k6UJbkM9osClCybOsnK17kWK8s9s4aSO+SvTymAla4oGM3hWgdSM4sPTIjePjOsC0Zb+vODPf0sD
WB9YIfT5oOKKb5dIBrdYIpwofbHJzyNIMf0C1h6e3ALFTYePfNdgf/v02SPG1LTO2De6sryKXhAA
LIAY1WFmzch7VHjPuzd0/vZAoHxKqL6WK37TFrnY7IW63bTCwXsFvtnJBt4DdrcHq89vSkHct50x
fOrIZNI1M144MoOxkrOiKC0OaHQYhMaCbz+2/h+S4qENAFiDhqBZ6kxK7Kl0wu4JW2L6+WIDGKbf
oSrumQkk04asCS2P7v6PBLdvk2g5tQ7Bk5StMr6dyN61eU1lK5GsZzFQmNCoE32X/jeen+kTvAUN
uLrBmrHQG4uYAFXymIW7TiUN5kw8RyTyQiE+utZ5tilK1J9XquEX6BeUpW7UTbHNzqFjFn/PA4Jh
wqhKj9+iLqR/89ZdCJe/35RLHNqWqoT+SKSURLBR/u0gtReU/u/hypXUm001lrm3SZCvL34Lkd7R
kdPJItkTdP/RLuseMMEvu35+4G6ew2kTLFO2Ir7KBSIkNk1HJDaed53JBW39Gryk/L0bo/Lx/6Qs
1uMwjjDDV52sDyt/lO+sjvmHICMn3bIxjCCovimIelE/P82kZFXjVphus9V+bj/iLibudWvDbqDB
kI8BeqKv8MxJJpnxQbKcvWEF0HXvuLdtmGAx5ZKMbWlPwTo7Fg1mGacchXqo6R7lEJO5fMg3A3mI
0Ir7t+O6+H4wdmgadtAQYfnaAQM9OWb229FSH+zuewZMJAI2NcXK9afsQmZx7uiD4DfsftTeRvM7
aCxUQh2RILrfrbdncS22yFNacagKP+bwsMnpwqm9x8BxFLF7KAmBoKO+E4vgekEV8nHJ1lJA2ZWF
omBBguh0uBNN9I6dJ4gz1sruA5fF1x/4Y1+acSLC/s25mf1LnAuv2YGBv/HkgLp3IMRxh1tbA9i9
4HN8lwQ2JMJX7X+Rp2SlqVyypSr1vZhIQZtBaO6OUHsaEvXz4lC81MKWSSwnVUsITuhaH2m0xtTd
4TrWPpuqFO1zijj3C10pelB3JB+ZEZrn6+Bkg6co27ndshzN/T+zZCMswXX1og6z7eMEdS8FXkxK
ELcOF60XyoxUV9zJxEkY6boax1tTzF2QvWCQH3QrhxB9QW79CUgdHWTg5ApQf+wO5VI+kNwHeyCE
NyPwTr+l2OqAmuggSs20QJeE6hOVhkl8T+q1SHuo9NVFzkZqQxrM0whioidjjSATNtLPL9jLUr65
5sh8WjdijufezBTfhTPUunFchsVO4p1EFFJ1CDElvCpdKcXl6JprhM6/XtugBE3+qCnqbjWutNHf
F82eqclJj3CgW6v2WX0mh/P0+C5tIl2TbCc8eOKNtxL6o/b7SOzMBa+PWEXGElQnauWLFnJEGu0w
EwdhUlb7aMz7+UDJhIs8x5rdYNQLK+LnVBNVcssZJREGupjeEzsC4zNC6opts6w5O2TvIm85+JdP
jFt28a6tt67chbkjFztMsbckCUek1qKShwkFrO8JhuRcYsbradD82BuwgTuDVZ0eb+zGsUdJpOE5
n4w9UTZ2E/NZdbWsuaq16uppeKOXo8GOyzZsn5frZg3jwQXQYSaQ/k2Xkjk7BwnWS3rj0EKvxRWN
3/SvHd7jeX74zV37AZ2OjMjZFB+BwAPIO2Cx2HDNaHZvQfvSiLG9UGn5BCE2ty6I/431qDrvhUqf
wSzXBlJhBOEu8kp3KV0/WFzcw2eyGrft0/NdORMUMUdFrwCBCKOazpDpyVKVE56vvUWCCjDxYyzd
OjjDoL/6zmxkoqmMM6/5E8TgEkQZhD118Wpc9csbaybudTT4bO8YsiT24xVsT33FHzdB05p3uP91
UxTv8TiwjteVc1h5Arzf5Q3FVmPJLgKwkPpIilo57q45DXfneyG+Dnf00D2yCM1MHCAjtQzfrMSe
vQN8oRRoEeGjIoKMGPDnAL/IBQuIJ7DpnfIPTOkmAAsBH39pfID2JIeXGXoi1O/4/nDQqbOhqvDE
dWFI/83ak5IczDNJPrwYeI1nq79bf5vZr/JWdUADmmbwh2H6viT7dnQ2WFPu3ZaITpPsoU4Sl4jw
xd7AufLCEWww6jAaKqarlgNxu6onhdFuTlOJqxgq6B5+uyg27NrArNTj85uBU7oXBQEESU5bNNAp
aFjI0RCE4a3Xx9+jXcARV1In8C7T9VccLlqswL443AfJYXkyWvOV1BbdOiUrnncToRwvcAbRtJ2Y
CnM+cjjC5Y5qlDJkU6e2I5CasL+jiOIPRoHOedbHwA9G1xE11sVDupHK3dCbyoW5poKYemzwZ0dG
bgeNArcuGUHTfJzu49hjSB1/0r9HcfaNVY862fBn8HgqyfbaFrD6B15TGd5v8TEnA72ybqqOFCmX
79OtfOhbOLl7Z5c4oK+Puno/VbMgq4D3gwwsGVQ8GkobSNg0jriUD1Gg63qDRiEplK6PPDKndmyg
JEAF4ur7szn3LrFZCg5898Q7TX+Y9XpPhH8OR8RuFx4f6EQFby+XGxFrvFUzTOYeDK3X1LO7XckD
N0X02J1wgvyOHdXwzEL9hBDx1EEsYcK6OuGqMY9ju01KU3oQ5pQ9ft+R1Oj9RObISZrSqU/DEwOS
eOOiANL26BscXWhzyAAtpHR8nupdLxjRhclduEaL1E9wbVzMQTMUYrGwDIOEXdroLc+R1VQbXp8x
PPlP/Qphquhu+WQzUSKnUi3/1RJV4rXl92G34fLjc4sHykMrixRI011JjR249MeZHztp/E7iob3b
lGrmatcqaxO747h5MKoqNoMSO1hQN22CkvOcULybHY7Q9hQGMB9SXJSWSZgwNOH8YV3V3G1+nLLY
sUd6Mka/aTkOU6nSZO6rLQZ1VMrXehHx4pJf+5VugD1ZZcYfu3ElcLtq+ipl09WoB6rSyHX6YYhF
1OYOQlHZwW2Kd0puQKyBWlNd3JwtpTeNhZ2tjlFvyPIcYyuQx29suyA70Z4QMhzhB/ZR6fPJiKGk
gKb+3b6JhhGu+9t6LvAEBt17dgU1KCOycyIC0DpBGICfZbl9rlpDNMEJcJn8zlzbErq3KRK3rkLQ
Kmc9GUFqEKo0gtnr/8RmEiG074xEc1yyrM9tUIKq9AjN7aWUs96IA1oCKVktvPPVOtDOjrD2m93/
U2VCwmmKQG4tCRLpWNd9+5PDwerS9gpqbAXM+QGlgVddLAc/V2MyINKKuVf+uH8dghZUQUxyLHY3
zRQ3uGEuwjxN6n/TnfMvVgIZmtdVvlOOwxDQN9kBARhVywTeiLrcG0qvaLuDyY2+xzwU+XJvZeSW
OJBq+DlHmMOcV6U7VAL0PQLLAQxXNd++4lXyb/1AKgV1+yoEUWwcvCNA3tKszJp8Ic1Ctcv0tzqZ
k5crDBxWTcSZMrxVpdEYVD5+XY6J9t3xOKSoIG4zayFZ7zKJACrA/XuVeYPAS4EBiV97xSzQR4+n
LrL4nP01zCu2ZG16ffJiWRPCzo7PsvsoL8fDpNb2qvp8RqLXL0MkTuy+yzUxt4/kkleSW3st6DNh
WZR+DHNmhWjTBtCCMBn6XCEN/SjBm9jBTIHSZJ0hstMwO3iWFjq/CEZ3njok3wrKPfvbbiSmQG0F
215RCX9RYKKCuhO+gdHa+muedMe+0c0BFOXu329MFTZqH/NYTjQxJuhVXw0/t33lA1TfUIc9gXo3
Q2G26UWaGH038uWeml3nYtpDW797ZBrgFCFycrcLp5oAG+LfTbWr7UvCGX2Ip+7iaDn+cdUp7/m1
KCnln+EtQmH1/JA2CyiDxlNLbx+Ma9UylAFE23NxwGQve1mGop3LD0PO5y0kCEU6AQBtCxtIQdCY
XTT6ahAEHaXxIgYb7S6sqWt6d+MZbUZ/hu34U9npOk9Zbsyl+qUekbN5cxQw8PvEt45Cgy5qvFUB
vdOpXrvAjmwVapU6DqHYrGqPPIDkbSTtZE50cUwIAeWSC3JnLahIAraBtXRj1FWGqBhatmknyRPh
tasbBZbqAvQzfaz7CYxuL5ciQTgQIT6TjdGB0zhqhTJnPMCJoi1F4BazikD/PQ24I00xuXTeVOTG
q7MhDlGJvP2hVmq5NZZ5w4MeoYXh1mAjNR8x/mFOBGq4jw1vv39Fy/0h1ErHd+29VduZKcyU9iYV
5sGClfTH8C7cb9c8JhLG0Kzhh6ugE+bJUuUh+UsYL9sMzUxD+Hr3wHgkfDyCCyRQOPIivMPrTJ8+
OomOqp1AJZWtBuqPo5K+k2oNTYxsIVnSAH2lL5sKyJ9agyAanlFtSbTxrPOfgTP6LcpyRayrfpSm
qd5pmXAvoQTWPdxLdP+QemkK5LWzkcF9vM6WzzXeojWvmWLIH/henczOjEMw8ZV/BCLVayhXDdr1
iFhmnVnwdB4BLTX8rCuQjtFW0FFNpbu4gX1NeJm+ayCRzJCPpa9DQVFlqrlMIxKN7Nr2goVJf4uI
vLiMHUh1gRByhzfP7iKuRS5lseVUSjOyP5uSsIzd3YnoHV1JNkd2o8ekkSKtwEKlAcUQOS4DGMZZ
dXdt4e6z2J6gGQBZMP9+lyyZA5Ja4C0ld0Z1uTUINFB537zoIhP2S/IBBUeOj264c/rfeRsoI8Um
bO4FUHrFp/zqnZR36KXSPslzS9m6gb9Ira55Km1N+GtsahiYhKa1saJTro18n2lBcCaTnc8hAnLY
D/rJVCrRi0TjLipnUUzTr/RWR2amxCKbBXY0lNdRrlnY78s66wJb6a2pTPlgR0ZgmN8WTYWmHzOT
so1Wxc3CIp7vnHJAytbsSGQg+Gp/p31Rk/X+ww5vg7vh8U4S2wNoONs+ecnj/sWXnsl9XfpXobVf
+47WjmjTeDKmUMg/1iq0ycM/7T1Jl/N59rQwhQmA+URXI+RC9EEb/lkuLMkTSUm4Vpdi5SojDbVU
AWEVvzTKpl8G7CbpNwbn/zHK0q+r/6E7/kpC26xFVzGQ6J/xyAQ0MS+q2wMamrAtqT2bRgXsY27J
cgwBm7vi/X82BwkmTcONo8XrtTbKFkQzKBYrprt1i04ME+EV6zxtIuaROYq3NCsGrPrStXH37nur
ZzkyAkop7e8P6rjglsXti50murxWiARJd19t5cxozp6EroR246PvFPiNAp/NmtF9wDefJb0cJfw+
/m+mBEaTiRJa27z0Uy8DEjlYQS/3o8WOQU7QviIJWTaYblySRCaoJbI4KKBMiUAiGgIQfNieqd9d
T+5rq4IXP6bmZXVvQDacmpBRIKlfs+HW2SlZvRuHYJUDB6Hm7XKR3oYF2IIBts89bl4ttf08r8pR
wvdp7LF7m6WWK/vC95uol90bGymoAVvX+Lgmo6RugNpEtswWzFnX5y2IVI6ZpXuc6wACmcXThbh7
m3/f+jeQyASCj9J1sMux4e29OalnKSMW+R3RzfRBkD/gNdjnJz8XBHlPfoXRQT5e5E9/cvI+b9q7
soqE8Vmcem4D89UlzhZtWIzKJW5qcff4eYx+3f045vMutkVW7xUXCCYaNqPy/akDnChtE5iNuLEM
258ppvInINYM1YM+5QhdpQ9ae2vFPy+fQXhSk2xFiiOsCUF5yCUGBe4GMdLe3EgCTtgu/I4B8jRR
CecRO0dvQgyLVmFL10qdAG2lmG1B1x2Gv3gGuC00azCwmeYjABqOTTqdbYad+7K+kKPNp9QY3B1O
ufim/bYtPjzy/NkxdBnqmL2K4KopvuSciABFMLFpbSlqwdBkl00a4DoguN3FfAI6Y10oRA1N2HFz
RyFK/O7z4JZ/0yq2DxG/+g8TL+HHRVNoJhOXADvZcXjmmimwl3uKocuKG+5pOJqfETfnfbVGXkt9
dKZFPkFg0WlPI+cphbdcrO6hwNEQr54VWl1dG//pfuAuSC+t46ui6VEXc6FOMJsZZjOhG8DRfxY8
yRsDnFvQGs7qGh7yU1Luf78zIG7lesg4Exj/IM8h8L9Kt3ZYzHWkdM0JuXhZENaQNlOIxXSaWLQO
VqR38j4L+L70yNPi5H4UZIvcEMeVPe4X0oGvE9GYuzMpFUPl5PtP7FJhVNrT1sAoYGXaqmauqaWK
MjyPh/io73jV+MJrxW0xa+YxOBFYYka3YIun26BORt3JZCy3yeUrp0f+4wJAtp8DpJVeM/d9uEOh
t8uB1jtL4x1Wbyo5f614uA3GSCCDwR56hyFk5/36TUAVG55K2YkbfdzaDNGsfKFvyNHGKCzkHnvZ
COu8rKAMGzxxz9erMcGCt9zjDQWwklhOr3B0p65pkY27xcAt6sSPEmj5Cx+OnCmdSHAzBfX1JERS
2h4AUiLUtjSiiqakxkoisG3GrXaKvjw83ZtHBxRkMGIvZMUK4VaxmhpDEvIpvzklfFwYbENIbY2C
Gsk7Mc3mb7nFwr8dQyinP4H7LuLot2PViUszrsWYSbNkFfqnqR8SGSDviKbD5FQ3ZfVRCGuZoH6H
hcnra/VAPIQbKSng5Kk4Bnk+srHt5q7659/K+tTkucHk7uDItTJ/IRX5jrYEazhKDAiMsX8Yyf29
bbbVNZWXEGPk4T5LYrWkwOkkX8nkGPiYQ6I3xzEZ1CxaFA0Jpz9ymJlQHu81KbMIuY5BsN8GCrWn
EL1R80ml/3pOShg/dYApFXMy9FoEBsgTKcXMRfcO+tA2y5lcypcaxfLap2eMmpLs7fLwa9GIkMDo
/+yUy3F6CHpGeLns5safiDZY4oLxY2qC/18ifSsxq87lsevD4kJGGl4enUdk7H+jgjP+ZDhtZ1bb
pDDGYGmblQu/2UBTpsVfc7OuHfKFpe7AmWDPUNFlaifju+ricr4NWxPQmedslDq7wAanDon8HdRZ
6NxL/EUcKqtsm25F50uhKFUHOVoslcpzDxyqsZDbgGd2NcQTjtb+TPAqUSfiAIe1U9bvKw4A5bLz
btliky4+6/JuZmLUDaK0QuFm8l/eg1CQxpybHbp8QbtZsEGvmFA9obd8eXF1BYRb23T9rMp+r4fe
RhkiEX4B+bR9C8yqOMZ4vVk1LRJdDeDZA6WCX12fihg5AYaUljJfPtWwacqrPgOioOqy6qSjCuyD
JdtcVNzCTR+NV9qEfuWpBCrO1Kt3OO1w1cuUmks9XQZFhVjBglPpCB2012lAxI7EqcU9JJWh6pko
wwYP4ELcdx0F7uzY7tZjNBeDZT1iOG09yJ7BZkZ4MN3dVNjwyeGkejWr70N4soYYlPuQ07GNX8px
vuFBZMDYwr4rE0YoHCvVLz9z2KXYI2rW0PjI08WMjMcW10zV0+ZekooCTK2Fnys0D8WWv9iqExou
LmOcIJAM/WiAtlUAl+7pyWoVxXh+Q+VeGa3nBHfGI652BqhGQogR6l2HUjY3JcpcyehVqbUgXbLZ
VjAWUGp8DCemreB/pw9B8ubF8ugiRWpdBl0ONn81f2w4jC1aI22+si3oe3k5OVDEfpZxzb8PSWo3
EToGHjuhKPr+LXNE6tiKKYDexJg61oOJnfJChkVJBGtCy/bTqHwhzRAVSqJ246VXTQiHnzB47Lz0
gsuEZJt1HnsgH+ATvFw/nizXxI7U6JlMKGoMXcnqLfXd6BKvVfkWXMjB+srAl1JwLtznSEypjM1Z
hk1pw7xR1e2OkG1GL93ZxGnpEcWkU3lAp5Trz62HZ0dXONXMIdp2StbkLDVX7yIrTLCSlFBUqQh3
0l+wrXDNTM5E4Pk2bAmoaNj/JSz01x7IMJRH0oVE2tZhfJor3wAtNlky8uuF0q0hl/VsYtkbtARu
+krTE+INj9G2xmF/+TaMhYotL1paD/oqq6qJ2OQ1EXviRmBFL194hjJFjwCZI22k1MgY1TNZUqyi
CfxCR0zTX7gQErI9883DO6zodFcTo3UVwzXMkXEvB14cNAXka1kU4FrplbbRdw3kmzfaquSP9iyC
9ec/9RdhYXDkcwAScCNzl1891m48OJmxMqgwqu3dooc58rddCoJSJihKRjRO346oMTcm3ZUOOVdF
TVBCryhSfuG8snMIUjBX5GxWmlWPs7Sw6qOYoEKRDeoeVqcXtdtcEXmL1BCBlFrPRn5foAxxUz7a
IQPX1al4kp8k0bwHL30YPf17PPvOamIeGOPvIQkPbGSUpU0mRpAFS3w37XRoRTqs9PN497tcqXru
bJY9Zx/AaE2Mld8yplN54suEAtAYtkr2tCNqfoASet5eQHJzsrjrG+39mFrzbYdMDyTcZ3WT+I0Q
sXs1lEjo8GCkPK1vNe1gUd2uj286zaQa2CTaj52SJkVcatbCPH6po2rZeRGpe0bzymSncRf3LA0c
aYYpZ5Ci5CuykOeCzcyQQJUFud2lv6bvsGAKujTeZ5cDqolpAVpMeFwby1X5HMKMchZkBKXyxz6B
G12/snwZFVKB0/tBCqU+sYvdyXVsyLsij2mbpmYo1bQpQjarxJlDNlrDu60bhVGtvgf/i0z2+01H
J0tM75Lu20hOcsah9JAmMA3IOKqGb89s7R7rzksMbeemJbv1gLXzgYdxrfsZuL1oJ5gfP3I5uALR
BYf3mSgq9OtiIPS6VHWv48vPv9hLpZs2dkK9fAKt7EvqRXQ4+/iLS60ktnWHntEhjrf55KxGDRMB
jOrFaq6sZKdF6NQ7pHU3yUQtI6D2exrQ8PxbXbztdJ9KOhJGlqHZjWz66ruZNAGyjmAj4hJMD2E6
j2liHdF/Z7PWiVBX9BcPn7GIvKz0jyaw0IYeahfBKBgMUA205glyPRW8lnriEb2eSd86j1DLPPrQ
uNNQR65rWlA1Al94CIlY3RPSuQMJ9WYlXXo4507QOHWqZaKOJRGpesGsW+AQBVU8j0DDRVKVf1o6
nzWnfDw5RqF/vhB7o2wLjw6ihysbFqsRJrIlK1ggm9APSZ4b1GRbuwACGtJm2GApdY1Oyl9RN2Z7
Rn7ydH6R16MDxaD4OedYxREgXKGprYI/zR1Oh3kvYLEvT4CvRfBbEfD6wCruVjcQD1UkV1bjCsJm
/+rrJl1ULQBzuDWR5wU57LtEG/MI+ZqtifOeb907pqFn+j0nKqtHuFB1nVA2f/8WPZf+MnZrYOxA
pYM6UTayRG12Q200Y3MWRRrRgfQTF+edp8mW95GwnHWlsItn3VjScKmNeIL0YodfFam+mJFpeEKP
eF/eq69PSMcLO5WGxZBHnF+I6pCCHq2Ja1L/hD8leObrLi2gWCsArYwF0PCnIsFBC8OOHEUYVH+g
uV+XUS6QsM5H39rU0M3045JyjPX/v2YTr0iZtK1jAwGAWo8f1ncRCF4L6IzK4LrfvBVqIVpHsRdo
ttm/1/UC7rO+DEuNnzi1T2ANV1e/NtgkcbxxsqUqjnKtvxzFC1atSbuFuv4lnKfieY0OfIVmMeGj
0ld8Em5zLelv/Nbmo/Eq3J5LTd6JnLehr5039qY/D550MrYd1EeKOmvHIJSayGTag4G58yqUzZww
TG5aJ1tBTN9pGouOSmZQK4Lspr4Dl3s1zkAq/L2ywCWFVWIQvhc1NotcSucY4W9+lKE2648FsBeI
sgRAq+zsZlZJDESuZSyXggjyLA4ZUYq+bRm86ppH9PsXPs7sWsvycerXx6xGBJXNiEyBUu2k5V4C
jxxAff85C7bdWIf7G4ETlqcmsmWT54QMRXLPXOS5/2vs8f6TS6xcG5vFIHtGNNKZVPS3pxJTDWnq
yj05uC3xzbSjuwUIfel02grIHel9w1DPyVCddWfwCWpJsSylOTyW/GT0UbdnPaOFjhmfot3F9Kze
7Bmg68XtuoGBiL7S6H5Cu8jSFGCA4v1eTzOna+8+Pm/WqUHLfU9lBRRMphZ23ia/dJdbIr1L4asp
DGBTiPuwE2tNSAWBUbnPOvSLF+HqMlFujE7DDtDDs5Gcw/x5WDMSLVu92mjxXOGuQKbs1F67BByy
1IYvRzIM7yVbJ/2qATxVN4tp3lo4d90cdFR1L2r4Z2xnJGfdeKKhJ18Ix+pz/3zm/JLUohe6bSI8
qwycV3fTR4beLO5uzP+Oe6jHqww6XTJC6TI+w4chlLIfrtW8KMcclrvbuu+OqtoaEx+nYGvaWyd2
nF63zMtiWKeHdvFloIBQhZfVUcSeZz7QbeWW6gh5hy8UIWsgs4MEiq1+VXmojXnxe5g7VBqlCI6g
iS7O4+vEcbK7yRuEH7Z/Rw9GWxwypHQxD7bsm9oUcNaC5CVUNORj7njQQ1A3uRFkG8F26vohz1HK
CtZdejsmyL4SMj6qHGmhfFG3QSNRUh1LGBsL0EbjnzxVKAbz8EH3APNjxqBc71Pa2ImLbDgGh7kL
OuYAGO65odPrb2bnTdZ5ZD2p4euRYELTWmKE9hvJt9KOcDGwrvriufcGFSnvgiNP3qcbw/CR9J20
oh2O5L77mnCzaAjppMt+iAvQSChyzM3+z1NFxBPfb9CVfDTvQIWha4NihdCMj0zLI70qTocGi2Te
7U3VnaAP1DtaKVSjzB9gXyguo9Iyfkx0Pv+K0VIw32Mww3+seFS7FxFeLFsLq7I7HfEllkJwmP0p
3Zmzi32c/bG7qy+K/RqyuIPPWp8JxMUNpko6M2cxZ0YPNeSbTaTNIEXUeVOyzHIu1a8xbJBqcaw0
hyhkKflo14rMDmvPR/l+SJu0ByaCM5MSmphHv3c42waNq6YOMTD+OaThb5rz+mpPl1LbaFDamSZr
XD0Wx6JioVc91pacISDZUCYgKy/zfpF+QS5ndruvikqTPb0t8leNKCSq/du4ZqUjfoqSIcPofqY1
KSdjGAFr7Zy7HG9y9WMgXeryq9xeRE9XuGN6GJcGzIzFio5RRCO8bSFtQ7PjqGRj4hYBvgwCaQH2
UsP7Ak6jHOa2lKPe20ilcvsI1sbp4soaG7ve2osfGARYyH1arJxwiBJTSNA4aQuDz4zm3kt5j4wC
qp979SWK3jaWL11LcAz42SeKxOCCwQqc28VIOWqc6cmnCxrHiXllrEE+uBdYtgSgSVcGG4u7tMHI
BelgRllqzZAWO1wwah+n2m+ge4WXITEjgfQWeGbhP6avnV8jHHJ8YzkJg8ds+chIjPvw4PqohFAG
58J3QC3e33DipQAzVXNBGzDE1vr+2hZ3Z3FxuiLciar9t7vinL4QkfoWESAAzw2h7nBsPxmjeZBr
bwt+pnXraZwEHNvsFZfBoEOUfXBrdRjxpfBY4yvgqGuoTZSw5ury/qRMhpzgLjh5GCJK3JI2V00Q
jlp94+vvnEZjNvP31Z6KZlK6+6pRmouQxAZuQIJFlv58Uf8oAop+nd6mYAdS0Uv15JeWKyEb+Zn2
oKnXqMcsvmZSVp1eZmtB0V0tEByS5EpjrjaIldHbZ/EW2+4ozyH27OWGbUjb0j6wunOLE9nRzqpj
Xhp759n4u8L9E2NnniMcrvLdb13Brt9It0YuL+O7HnlBoKE3MQTP1u/BLsYs+Y2oWRNoFTLxFq+X
/GRuddsnH/ndn1zW3S2c91t04vPBzKvSq6AbCjuRLx9nwnW+oAUiKLhCrlSV0hbJcnmH9n1EbUxn
w6cs0Oh7rk0VqAKpF0xKpAZ9NtktinJjAVlNL2ipluvA3LLP4vIPbIS9jq8lCGT/baQ5yzyiDzTC
r9LhGwLRpE0/pq183C/QuHhP/kIykytt8m6+umC6mRjxcLAjEKspwlubvU1luAkWQMvPnqwQ5scy
NzYyN9j9QqY7/NSEbW/uMGXqw3eVpGUKOWNL/CFZ2dfHJxgdGzcWUnxxPo/FDJ3pHkdm/gMSLwqH
L1APw3hq8H4CisNq6dBRgIf/lMp2BShljZEnbI2BSvuixVoYZOK0OzsKUwS/N4pJrO9i2WmnqukR
ggJ22sajRGWGrQLWUlAFSOpF7xbznu4yVO4DKmcItFwfIYEy11GD4E/aWeApVTTznljR6+2wweW9
YbAeSbNWoGudygmZ7i7OUF8qNQYd6rKFF3gb8Q2S3lXoAEXAE8SmK394ADPP965bbgqRtbfSYPt1
GDz+C2H9um3gIcR9ioMDX9N1yzXw5XMylZP1VcbtEVQoCBGjaXMCylWXfeh5AnPecAFCLnjBr8Lh
nM2w4ikIf6GbdZ233UDN3034MFbNbIjj6bAFzms8u66GQEjQ7JxBgSvJAo9MyFXiCYGsQpzw1XN2
wZvnnD8SZe2uJXtjDzQdjjghM3jds76YqmrzJhl8rM+lfyhwHGkSo/AQ4qyIqdldNfZ6IVUIXfqf
awROf9EmWjyeLiECDVLBVM1qCgSFXFJoBBYS0WeZ2HRtavh01SAywlnx/F6D1QnTi5cqdc2DVIwl
fCIwiquYckMzmCzRYXtAeLqbpMPCWFEEuIe8iJL6SkBomIM/l1QhG0GONDNGLRJeKLbkVU1Xh2vx
OEZz5KdE/xqm400xtpLFOqhSTHxL9/epEfxifAH+01yiPLTuLROXAvQiyKuTHTHfio90pfT9cp1u
KR9Dw2y/LNryz59YMgMN6y/QyMPVt0IG72AlRFMyzatBkfGkvBi7X2blq68BrarLQ/boKaH/a9Py
uUQy5cG2b8n6ZZzDb/vEIdVeGrkDqXGSVvth+uk43w3W3vHZIZ8goHHu4I1yFOfLilW/iC9yackH
RCuOOc2hhDg0QiabAhhEvXUp4QWsMfM54wUXxC2iLi7zLYuz7od3a3f4Ubvz8zXdqOeWDmqrcTP1
u5Axc1yevbmPgkOl+qWTVVpGr57gSdkdG4DMFDJWMaVDDqFJ4F6p1I4sve4VIYykySO3NP8MpuJH
/116lNq+1K2/fU2+z2FEVIDNZHIb+YsU4PmhLb6KxXw/EoHXh/Zxdzc46RZcHPgaVmemCrv/OxIR
o3TEqDx+wvp61t7jLbknqIulNRvzwqIMahSUD1hrDAEZpm/5eVJk5AJnCYovwglnLc9QTLemEBPa
7l2AlxcDjLi2i3fIzv0g1rg6VD5k4vi/CF7zj/y/vD+L5+aiJiL5mQUgcWd40ZhicVb2NfCjsG21
H5DxwX7SC0AJhgrxgWMKJHgaeXuNt12igQUo4s4G6QBr24d5tf3FEhLcvh1VGPin8W8K7XVCt8Bm
22Wz+yyZ6ALpTEGxRIaXiy9cj6HkWclopLM5U9u6R1uREUy1hPS9WvFSQLV5bsUNVcc0+dT/c9b7
GTQNgEuijdbTDH/V/EASy6qHOxlEkRtlldYS0t0XmJ2PdpiRoAQ40Awc9YUkPgXd1NiOvEt63vvn
wziIEaJ4bD0l0tzMHnXsDEJ+/ST31Fiz50FDzq1Xs/hdhPWeSvPONyoqW0Io4nPSDxx0Ehjuh/rU
FsRSIhpV6r0RdZFp5/2a9pWJK9zPN4oZ5K7Kgw9ZmcLqboASxAgz9y9F9DxIKQpqelxjF//48Hbd
J8hweN6hKtahAWh2eqR2QezTNe52/4GpLcwdHBqeCROTyFF5mrBN+7RgkD+CUXwZVAeegtGc2rJF
9ha5X4j07tuiiCG7sYQRTQ/FScKWEwVm85Prbu7K0BM/0hHZvDq6NoNUn1XuE04o5HFJDhCS5WDa
qTxLOXYFTwvy9/qYp2GCSlJQDPSFNFnp6RuaKaohaWpB5eTtbCWA8bcUDnOvsTs4/LlVqoFXbYTd
0fIyiwpQDswnXI0ezrXP3gIA4LAYMHn8tyxjQGJJLwdllY/+dEwQq2v+PkitJoNLbuZfrAvgBO2F
1Mj7OvyIm3QMGjWhJTdVcMV8/C1n+mBbTsWzWosR8wNdSOHH+x8qfcOg1NPAiQPzIUdaaGt5OOS+
EMEQH4FXpXDs4nbFz1Wt6nWEjF44bQUUukGZY8FXSEKHeQPNb9ujRsmfClUMDDoBjm5niFN99weT
BWtQQvYVnCIXbwJL/GYXISxSak5kp6LnRComDl7BHGrkRmf8mrzoH5UYdBbS4OnxphhZlTCW5DZs
aDDfkRxIKYcxFeudlF1oukAqNOIeAp8PI1ToIHtXGSx/U24nYruAdUCN0E2iTzM1Vff6hS0yxgfP
qjjBljQAi0W/4+ChJ9SjI9b6NQh2PXBCdVSTTfhe7zEAs3fYHmpXlByedTwvAP3U6/wmuyBBcKMw
pPB8/2eYaEa1D+M4/L8chl52jT9SPsS37L5T9mgvmnC9cYKDZJ0fpAjbd1fgbBPSAbKq/0kayEXB
MCLQk7lRyYoONko0wGm3CX8NmwuWIuGnujVpZ71jqsZOjINJVlrX4BhAvFd6m9vZdP0t9mWv54+B
aL6INQ9yGghCDIAEBQvxcRewSxZHGmW9y2FJTvLxEXNRrZkbnGPxznQ5I68mWuYY2o4GPGxhoeTs
wov5WvftJ6+atSTMh5hxhpFvL0tPEIhkODpJM/4RtR1PqOUwN/ZOyDhkFCtFBptdYKxa7p0Af8Ag
6NvwS58hw2gPIUaxw0C9GKFiNwWMabvv+xg9ZenDVXO4tNryqPBsPtCjFWR2WIHkyzSYeQHiR+XA
OOlfyziDE94W+WY/0cDQWtkYzKBzGTa/uwth+azP5lheZOmOdd/c8DQ35kaA1lMqQu4+YdF3Wkh1
Bxvatd1lXZvri9H06dzTv0XJCXnC1gwpcLT2AZsNe9b/QKEj97DwWqDjAK0+wJzpEpoFU4Ie9mHr
9OykXMY8u+OEmLIG5Eue4wj7fWXMwXKvjf6A7AAYnUgukXApdZSX1Wz5GMKYiOCUZc1ae+n1w7q6
hjeSeDImIM+69VUNq4ZBNpP0065GT9rlgBF3wW/SzmkmdNEd15J+N+W+szHIsYeJbF2W9uTGAA7V
sYpvwvualImQNJ/0PINKFYPtjflcj5UPels4OHzihL2hU6IWbPhstikKDUAUSNA7gaiHUdUmJh03
UotzNv+uRcLZksDSS2NEob+B5+wCqGEGeEdkLktR8yStElkYywzaxRUZJCxKU7EgdWEZVkIGNB/0
mTLjUA8rDXUXZ2yxEqz84zk9lsf1xtwfHfgUYFHnVl1Z9Hzjhoy0mxeSHPRup7ANztmmFxX1w3PT
FNKsQI1M2UDJW5WErod1BgKeMCFqRzjTbHTDbisHY2SZtItYkIlBWnpTuoOp5a4eDEc1fZbM6DJj
jHJlHel8iQ0fpB0TBPspp/Xq/MYUHGngHBmxyj1XiwHrAfQCG6QZIMlVksH8ikMuTIAPN6x6j0Ib
Dk++yXA/1/L/ooTmoaVvSUXHijnI7DrYJmJEDLDD0ekMUIF4OGWZnHfA41V0AupnThLHUakTaOAA
897s9om6B2N7FEwyJpRbc1OKZAD8Dnb6ecrSxsUV//ba643X9ABchyAXzuch5ial4EQv+tZeNENM
/rO41PNM0M7yOsUpKwd7xihaGbMGkAvjiSzo9EUgZ8GcuE8W/cluyBowTIpono09/FZ9ooKwg31r
moTJxYEyF70d777JU8FmmusC7vO9yzUQoyLGvRJLZJApHkAsBZmqbHbDuQMWw3azbXxGFxxRMAZw
wNhocHLt5x3DdSKSMOKmo9ZcH5OCAmnOP722EUAqSfNX1G3YJdWQUZUit9vBmZOePmBdgbpy1d0W
+R0c9aK4Yt6BFzaX49njNwEWXzK44XuMW6cBg8Bg/rZ61i56idS6EaaTUu9b+8Tb0y48AfSRcvaN
DAiiT4n6rmmWTcr2Iv4qJe90QK3JuhqdA45Nx7VaSa4hA+aTlbdo+2Sa+RsSGHzM2igcAJtxaK6h
Y3uuSuij85w+F6nJc/Rf9hj/OhyGwGLyhISZVHFE1gM3QC5b0HCqw6uVCB8TIiKknEOrsFQjtNOg
jU4YmEslkIIAOr7qjhdYHYdlm7ow3t1Jcp15xPz++1qvvdkXCdObAfIpWvhxMlXcaqjr8QeZAdXB
ZJXjbS88NdNFJdsXiF/xG8upU+DFCzIXSYEIVFdb3gW3O3tCRz4nhttGYutRXRcnVpjaZ7JdcPzn
8nkzOzy1e2lKAXNIYLyYZSYPhVVdoIYLXpIAKNdAM9kd+MS29NXascv0eMViHkxMlTxkwClaA6uJ
J9Xn91eluhnH98L+ILBZH+yBzSMXNpFco70p/w3/uPXSMeF+/unsYB+riy90aUIhIB9QG6GFgSV1
SBcMG6ZnNeWlYhge7kIyjsG4sBlK5JMajYtqThAYz2FLvXXQTARKlylHyv23m/h2bYQ8cHVwKc7D
56W/WJR7GXeOt2oZinj4qzISvjbtR0+KjiBkqNVBd6JnpQO5UCC2Qo6yJFioK9bvIQujvqocV9dI
xWPEa2IC5Uojf1JmyLQQBwd4L+BCITGw28BrQgNWko7fwOZBLELjyB//ZpUhLQTVNeftNQK5d9/Z
jknz5e/sROVclItqmdkxLN1+jIvvFlz7AbxRETXYpFqVbamPHZ5yI7Iyums3QHrQMCH+9EbXWj4L
Dzc3PhCVugV//s4NCYvABRZiZegIQPqNQJkAJsgafJdHT2nl39kO8ZGsvKBKTgxtn2Hqi/ehMCS5
6oWPBvaXpqvwAV1lSsgQsuuIDo2b0M8CMTL1ZfLGbepNNn0DFnUgPl1Qs5hyOOoVzPS9RJrjx0gY
ro1D0lJE8A9rta8S1eT53t+KiLfUV9sMpTDR7LLd3R+Yvq8cwHNg1keV1tfKP5aw/8z2ExtZPmUx
Kcg7YSHjuSbuoclmHsfZGy2PIwS4u8C54XAy/jZvcIlb0khydpltM8YN+F35mav54IYrjHhZz5l2
JvReg8v9q/OW5NocBDol9MHHMt73M6pcd0n0q3bepGzDKglarjRTef6sb5ixE2CFjii0NB3injQc
HnN8RFFHb7wrfq0mnS5lZeTJwtOqxOWdSzXNIGjl+65/wXZKX+bjNOy3XK77lR7kuuNuHBa3Sk6S
ecZ2EGyJxckw4XxyasMuXY2ZqZJL+hDfmJiSfFmj99IF2Rt0jovuivEtH7oxgQTJgQGtgNlcpmR4
G7Es+G/e5gchqmwEaCyxseWAO3ZerBlh4aEUcOzCsge+yDeoNUoxKtFnt6GZ+shfUf24LXPyLxmw
z/3CYwFwgodBabTv4ZSmEq5QEBoPyD6xHGpEWH70mS9COfU2y97rnJPIre5F292L0pGcaUiuXhpF
PGtYdDTfMFl1h7/Jo5WcCIg8c5B4oaNg+WTFBjTdhG/wsDXuR9keR62mtqvW0hh+IX8TOduch72P
OX7VBc+168LOYqD18R8UtkQuB0gpV6AA+8lQW63j5usxWflBZ6BuxSmno4wEJuOg7nuC7ZjkZROd
erIiR5ohYEqrAZUC5yESHGmOugUDg1/VvcTJpSRjELFNy8XiwYPxf0jmID8q7H/wZXgtIM2yyN4h
a+MLLsKz7bt7GCmdUoyFgdLaqLUl3tOyLXUMThF0JxWpM7aZMGEqzDHoOp6aOw9EKP+4bWMI2FJ8
8OG3JeLVJb3voXjGmwtr1jx2Ct729CS/u1ohmNM2FdUgP/clfRNGC2JhhmcEITdeNApaqDw1t/Fc
3fQnDPGzIn8F8DVLX+RkqdUcmOC2LJfgsAtLXkSnZSdYyIW/68BhI0CnScdNGnoN2QID1z5sm2w4
3GR0VHnCZAB1SiozgMF+Ve7jNob14EnM6ftUiNljWCBv70SjxwoAuN+iJPYex0yl3T9do774Zgjh
hXfkrz4fR/cN2arfzdAH3uXWuCucUkfwrGkFqgXsXhaHTvAH3tCLqKgCkqzyYXrEj5zntlkUTuKv
H3bwgIohoqm8hHmf1/T0HlEUQk4qb44ZXugc2TFqNWh0uV11u1LN7gyeeB+mrOVlwH6puUkA8tN/
qNOVS0Z73YmKY5xqbwfOTIWLVfbuZsQC+kE5+cKqCd8nOyWIOBdPtgtHvtnTKsziH9NJtEWZAF//
ksmdMjOrEiDbL228O4gjwbYkeMz7ctFXvmeJtjwfbpaU6tuyra/2xlPqiV/Jv8oUdOeARoO9zneJ
IE7V6SaFPTmwNafiYhWqQzaa29StyxDW+DrnJv5sYzVqBtvefkrIT3XFlYKCu81AIV58HhqSrAVZ
j5fNNAjsWk+1Ty+WjhCoMrzA63YcaT9HxNLgGFMtScOvQwWCyMzd820cY87rsHtCRjLdt94Y9LH8
DrOlX67GQZ5NIqeJaMSbNI3+RqQYLeZqMlhAU3c9ZNCKVDjrXeY/nA5nD52TozFxyaVKkUcW7J99
cdH+GKieQS2AMqn0M1xUc7Tj8kUgdX8AjAiuHGZnrC0jc13eYS+l5QVC6eEnmp9maR3u0U2VqxyU
YM8cBR8FOO4NgmV1sZEYVf3UsWWoQSkKUiZoxpVX9SopIe8r2RLqC8x3V2aoSZ6QKQT5RiwyOvd5
vojHzLezY/TtbXCxQGTll3qZHZL2LzNkqONZe+crUr5NuTw7CPQRmN6tOLELMowgMrvXDjZ77GHM
VGIX+kDxJaLmisD8kYYH7XvcZIXZDllgLd2CaFyEjb0rfwvqfZql++ADTQi2nXxuJextNz/KaC1n
BY++TPqPl74DZEyrCyq+4WjJxG6IdX624B9OF2xrLNlIO7UZtPfjLTW/W8vYhpsfy+O/lRU+K424
WAVwMMnTtMZeU/3i65Ocf0+5Hx34UGa++EEZjA6ZFuvuzBIScm7JCUrXdBF5dR/vwoQqQ4WiNR1C
432+gajRehIUOP37cYXV4TK7tP+cugY3v0TxY27HxpHN9Rz2R+bvIJt/qqFpAe39Y/M+RyYu/FaU
gJf224wWyro8id1F+oWyRNBTFRiJEean8E3SGdQgRdHhqcZn38Bsj34aFVAGAqwCoZRNnemPvnET
sL3DAUT7DguzneZMXgeX19+s7Zx93V32A4zdy2RWBL0HA0LFaI7Idtlf2qW1yE+YkElXeYoPslDs
1wKsTvD+yG+3ceoqdHgAKW8iCG9ykI+sX8QrlyrnL136kalikuPJHpkgD6NT+Tb8uTT91sqJNdeW
nH3klUqeWp68sKFobYtAfhK971c6AM5D5OvyCwgYAAeGPg7qJemUbx2x+Y8v2T0FLvKbeeR1/D83
ocw4JRPCYv0DmI0tfnaYuS6WH2qrXgKrYSPEcYXrDcZXcGO1vP5sjydlGdHx0JlSIzngRLkcRXTd
QbGGuqlDccXaRjhqb7rmIjg/h/twA/jhgLEm5vNTRmtxJ99aB/6QEy9ZcPGi+FQqdo7MJkSoi/1Y
E6wXF7jLPhCbMHbkvEZAYspT39+BZzm8JSz6fQpBxHXhEb/P9sAPsz/WaqozOBV3pjyBpixm/z13
t6IJMCbes+6lf436Z80o+HVgejoSdst47eYo1n51aJH22Rd2YP9XyKQd42PKvN5BMFm6O/CL5wrQ
c36bx8blQqasghZzePC4jQsqomvW9GMKmAbjCUpVaDXpSStX38VjcDhEnOEXH7yd2Lj0QFdAxRiq
waWATrqiokOI2+EMbcVn8NBF4BNEQo3qTed4Oba7hu9i7fDuowJ5XzQP876PaqOcBFFTA6Sh78ST
XV0bj38QWZ+8KTo77WVQ/2BqpO+rfbJB6wcjziJQfRm99dbkmwMlIdIzlxJzklnRC54iMxUyrmYS
JTdWOMVMB/87EQLXoBlFkz21ThvgtzfI/0K6N35VdUIm/m0TD33aJg2ht5qd9X0bzFUKSqDBMD11
nFgsiEOp9K/fPISeRBcYK5rXJDque30u9hNRAqOUSGm5A+OD+p2TTxwfKh5S2l/OKVOigEWdOZbf
WjrzhcmqSd9pfpXWlKDKUImEnQ2yk16LpBut6RN5Lp3jdGH2rM4lzNIJ3j82W7yZ+8R1wCeBuhYP
tW5E05Tc8gkfU146UNaTX3jz/beSpnOv6vT/sp55lCtriwpp5BeuOIToWwYCdwpVo3Uun2djEvDO
jc8ygTrK8vm0RoJXr9pCzIN/Vs8oXlXGNlLeQDpY2fUSvQGn48nK08MogJfS6wSCRc3OVIjJL7hU
5PrYsc2H8pUPA01FncK4MRtTc6YlRPuJPu/+J5IGcleFYKQiSSQFcdaccDD8dGH7V/FOsPoi8hB+
qrIKOiTZf+neidqEqPzMZsZreoQUYel24Dm0uMFygSaxdeKNBvze1zwDAkp9hsFxxq/g51tzKjSZ
E9HZ9qAcKZ9CQkl+zY91PD1Zyv+Q7tIeP7slctxIUBucBPK4sEfzYuMWc+2ukv9S8sm6/W81Jk+8
guJ04BQIPn1nKU4M3A7cGdW9U/PAOJwL0TwzWVo1+Fa7m2PcGGHrPnfvXwfLLyoSEp9cb5ddyJye
4cD8CJZKlQNGGS8O0496VeJ6bdkYn3KQF1yTFLbb1MIUqaW6mku+jhT0uXMbb+HH2E+blykpUFS7
2j9Gxl18MZ/aNYQgOGpo2D9Ms8n/cpC/0zf3ePGluGlBlq1dEwJL1x+KfMJ8O0U6WgmOsRDaxTGj
M/GkGp2U7eTKf01xA6x4XqifIiNWaeS1VHwvJVX3HxwOkBCaN59fv/WV9eXX8pHlvZxDnEgFA9fj
HP3VYot0KgDWblpHS/hEZ9hu6iHkAs+sKNjqFaS7RlZUdN9ZHdLp23+hG8QERcyMSb+ihWswX6Id
u0xhgkAjcN4Ww1mOoWY1ZsRB4GOr5uMaXn3dDrdI+Q6VreiOSkZQjFNxfuUPtcygO5gr1YemDMy3
dsu54J8VSI8d3Gjle/ttEecoFx+mmfGL8mlvFQvTSSvq5o8i5LakVekvnKpEE+yUYcTijyVFTy+9
a/rk6lutl1A6Uak/Cm8vdAanIJe1hfQz3oJzGePnfpmeJb+rxi8MshoaU0fvKFaI9TYuQRlbeQNK
v87SNsJ7ytN2c4iBoOs+QBFdhP+3xOZpWd1u0wDvIY7lRNZEM3vZmG8gQ0DW/QnycpZEYdQuEdpI
2SXKpaWqqclbRbr89dPiXr6Ln9+rL2vFcWjdqLpjltLuaRVB9Gei9c7c1pQrwKxCp3YIoJ3gjI2t
x3vIB3zn8M+ZlKZ3634nGwA5x3ohsbHXup3FsKxE4aJtAK+/Gj22bWrPOl2VVviM5CAnMCgGNbdZ
uhBiAe/sw+TiKfIijkfoqr1SqyOXBp8jHRFliLjb+fqhRT3oh7kZcwQilRY0Mg/TrodCochLCm3m
noMyXzkq7JlcdYUbu9t3az2A6N/vg2PS+R8JqB7NFcKLPlNx+yek6c2SmAhphKn83MWiZ9HdewP6
azGTzkO3lwXVtoz/ULlROnKjs38KNMCBZ8XM7kf4N4Z5gVMJFdfEE+HSj57DmX7NTabLCz3LKgBY
3ovVLP370XeKzOlieiMC19P1Kg9Inj5msqNLbDwnScUPkrNmsYgVAbBbZbzrYSFzUnmf2ZfQS9Ho
UPvphcozS7TLmWmxbiBHZMgHgZs5ZXpGbDS0JI5qikQeh9L7U5FoAsZZsSSdciuPc0Xk5kcfDKbz
T1N5gCsW0uxQa8aJRo/ecSYD13p9rzjnmbXw4h7cj7JQCfqzqMKPJbTqjxpR+w+sTVFd62BjTT9L
Qd7kvc36qGvfRLDf05TuzC/G/6kadI8nNtHrgGGu6qbbI/Yg+Pf9qpH9uZpoJc0mnF9+R7sgJEP8
X4+N5pFS2dAwcoZYkotCAla+0yRkGK+TJiTKKTmn1dh8TKZhQPAAV6FB2ovH11R5fEuf/lmdlbVv
HVoNXA8LdK9YwYGqr6TVPP5zz+wFnsCdDP0sAEWTKBDCGzlFz6ZBrXCxOE7PT8ZHml/rp3rXBa3I
QJmSC7+SrFpn2WqBOuwZwGM7vbJnL1NEavKeN5AadytCw31qnarVgGTSY/CU9NWAut7RdY95pr7e
K25IA2F7SAzaCIQirTjYM2SD83NUAFuXhKHZi9MWN0tMxUfj1nVBSc5Fjpemon+jeHLBw9Sabpfp
kOE7IlWFz+4/fV+TQ72intxN0RANRnMzDdiBpo+lpmTvG2mWlDmp4cgpK68BOFPMkrMy1EDpKKva
eJ/w3Pbh0l+ZZWoYFSn3UF5v3xEBLu6nu3VD+mqifCtMSLy5jElklcwJhbZve7u9+m2LVcDDqrAp
iwUekKde2b6YBWdhkV+7zLc7epF0EFdQsRzijFhwadSf+8y3hqMa/svKTIZHADEMZGsrR+hx/eIy
fNHOTvIbFT8boNigwMdB9sRlW4JWd2fWoipA5jF5cVB0Tbq3+II/cE8Ee4xs9H1ObLwdVSVI+59u
PiQuLiHiDUFiO2UHZF8yQ17GTamnrrD/1EMMaHVGM4FPpumwYHKaavxNOJsTZGeHyIaSIliYWXac
G+RE9IbA5N6Ivq1MVmLGXrK7D3pXp9xo90vTC1Uvcz7/jS1rQxSOI9eYibdSxJXXjL7fUtNCbobx
eDFyqtDh+0v0EL1ygZ6dOLXTtllyGjOm+hvgIrKSM6FAQAS4b7sVFb9+DrBE3cgYIxoZEzZHvkdD
JfISPOOSGWcpFM2KtKHKsd2L5l3uCY3a8c6m79bqiL/ExRA6ePpb1Qr6QFXK932tikRMkPu5vWmT
DsU5DTGvHUTp0yPM8tKpL0Q++KGX8dEfglSHUI4wWHY6Vc4habqQ62qQeT1AEwKY6AU9jBZHBdSI
zvB6nXM0B8q2zEuoQvYfVhItgEhQwmqrW513viIA0isFXYdPxo6sJ3f+PsobqyHnKVrrMj1geQwv
i3doy6PdSpUyphFm7cNUCWZRQ3vcyrreqhAXJh1tMJTlblBy6RUbLwnJj/W/VeR9hvoVD3AbVCJC
2a3nU1CngZxPwbU6rPSBR4E+OvXlZfygNMUj2HAHpaE4Y+vzS7mETv6XZeg8CvmSQ+lyLz2SFm3c
tyZVsLe9ZomZwECsK3uLTJqfGPaJiCzdh6tNiN2VHDvp8rZWPpGI0KX2dlbWIFfDLMXtfPLKcSdO
Tu46Mj+5R0LaLJYRRmnGhdNyxq4l/6zxIp6gRgvuS6/ofR8kDu1BFyTmuxfC0tuLt/LM8WM+VYdi
0EF1QygPUcbszIemVTWLwVd7dUGvwic5s7kj0tNsvDHpDppClTMA7vElo9Hi0B9Zo6PN985KBXEG
oGVU/CFYiZko7NEN0UcuJPrv+r9IxercUESaQSFT7nC5barr5oF6KmFmpo7XLzmKifGmklrDT7r+
TN7jWxnvG8EhvBKG8+i/7nyR2tGLG8/NXv7TZKiBYwdEh8y4/ePXvs785FNwYlkQRzwXmQRqyUu6
rsP5QyiW+c+Qn+yW/PEuS4QsBYImamnuZEHGR+PRgLPhdac0gPjccCNStEsyBoZpQj8mr4uV/uNn
/7faOwRXHAO+9bRqLl3pMpbQ1pV6s7UGcMfRZg6hnLTQ7qDRuLS0Wi+9VDouJZr8XRdqvN3WU3+U
9JnKAh50y1Q3wUsYb831rLB4rl4fnkgdx3u20CiA05vwMhOASt91XkRI1YcyPPVJ4Tq4WOf+WvSU
uE/ddIvX1+DKpO4vA3UdUwM1RW9pGTruJqVe8Q5DWM9jTFt2ZjmUsy4R1Y2fn2CsZs6cajT7GmI8
JDT1AthVZHH2GZ4AVIDVTjWTHckZ17d4ln73S7qYB4KF++w77xUJKQsiboJB7828rHwNw5uUIzcv
tWRR75nXMTOowV6K52N9u3dZ1m4IveFnCQIxKBlDY68Znfej4o7+nwAnY7M/EdEEthg2jCtXfV8r
Gg5n0SR5dTJ6a+nydgwK1yYlgaNiRGHAigruAOiV8pKE7ENQ7b1O250bNn32wjODWNtJDo25gBOf
j+BVRg2AaTg0StE6wZiKbv8UrYPEgmAV52gUxMe8MxrvAopD66X4inB3qE+brJGHrfRwpIykSgQJ
1D7/9bDdDQsgEq/pBekVwW6O0nZqW5UlaW/8cap+T7aa6H7ZeVZtEz4uyc/ZnBand67ZxSHQptZ+
wXhBVajD5fN3H5s3RDT+Gw2XOPkH/9ZBothgN3Lks6YwVHrxFBBbas1k4JlmVXwXw8dC2Q3RhA9d
+QdzYdpXzypia03VNM7iWr8rCAez+HQVRTzr3kwdQkRWEM/wxk7Dj9azp61BWeDvWu00BlUh4zo7
JSQspJbxVE2STRBedGwD/amVMFSZFa6UHlBNIcrJFf8fljgEG3lLJTHzGxIJm+JMYd/vSkg6Mqir
aFfWuoGXVgp3fY71UOsCBkjimyuU5XWlY4EFe2vjUcvzVlJ96gioDQfs5ZkCJX7c4pOt7FUscaqU
VqI4Q2mrpxNg5ZM3TOSOH75atEHAWO2g14DJiSUs0hnY9AuPK7G3qziuhz3zAVkS7gJV2NQdLDLK
PVL4AAXWkQWFG7xYMYlpctUq6jYB4k5FtBhW6EoPSqGuI2lEMpE1dPOg0vUSkr/MVslYT3sihg0R
vkJgOpLsfUBHnjWFg/SSKmCfv2V4Mo9T1PIsJNzfx6qxwnb76n45j8VdzZCiF9urY2Cp73xKWq9V
QpDBWEwwsHLkpyv+RfKJa76sWpMYJsriuG6nluR2XmL3ZZ59ktZwiZpIwDmhwX6dxx26kQugTdG8
iaGChoi/VD15Bh0jXI1ZpfHezctLaOgx3PmMPNQKBuKy8m/Yy1/QOCor/91jcKccGkHgJxhQPpR6
Se6vtquOpoyJc512blRIl9Q9Pv8hcEllazpzk2Z+3rONTMj5cY+WLsZVefkYzCxWHl9vOX+2XKs+
X/hKFbW6tGvD8kl/zhJNNCjHaGjzzZ5qGWv51FKG54HRXyFgT6Q6V2rW5rfKlKVjZKykKhFY/SN1
ngpTSkm2f0sLOKfByFDwz1qdRHHQ4CDxTqGftP3CvNEkjlzbpqlOrLB5GbAQe6xOLow9EbHFCJuV
0x6r1xZAyEUiqDnw49zQIoA6B6vyWzEmhjAko9/TvFKCOWTS0DybUTkQvHvr6r6MHQeZs+WmVVWz
MdV8bB1FmPflvWt3jThCWoYMionYFe8EQwRVQJyCocjYC6sagwcZbxtjqFBnNJECsTzjtBgAX6L4
Cc6M0ABXU7kj3ipCAZb73Glxl5vcBVrNDeMztS4rLwDdCRwfDqOYbeboX2txpG84IXxg1j/ViZfJ
tcKGxlpZ7kqDY28/qZnhY5d070+DDer8S3m1S6j9n1MgAcYu6xYSOoxNZvLd8gR4GhUxAXC8JuPD
aPXTVeAlmIV1+N/+m/Qrjl4qWPBkqui/ZDBmHJlWUFRhXvXSihBu9FUE4eDnzr4X+l6LilRJK5BL
vrlA1xeaj+HpGlV2sXDq4dyDBF4TvSbX7aBoZeDJbMJY3nXNBQVDNxO2ivQGKNAS6FPaMbKc+BJ9
ltFxTHrUMO729zliQh7/wt2JJYJtbxzJVJO9RV3X5xz3C6lEbZJ+Cb24UTXiGQ9KfJ14nCrTdfxC
S4ShPIHCWlEhCw0yPuZ2ZlYe8+28bP4L3pJOAKIOePyiD87cKY9/4uF84wKshrXPLfS4UONQByLG
yZQndzOwgixyv8dMkxFb7ghkeOOIs4ge7p0RuXGe/gXTIeARTZSyc6cNlZqf5sGwSYUjYM2ADUZ5
xrxh2SBzCLlzp+HbPfGxmUoMNU/MouwdbTOsxMFNblvijq4WiXCA1abNIeSdMnlO5H0AG9pATOb3
6Zp9rcZUioCPdNRU5YrlexwDelY6YPfAAf23hovseeHWHYfYyX11y+F4KMwKeYhGfYAJMe0lZxDK
06RmllXXzc0dKhMAUyzjTAi5OyKqfrMGoN0iJHy7xdRjM1OR73KUnqzjSwu73G9z/dyWtrBf51+J
z7pxa+z3snaVDNy1XmXcQhQS7uipT/ebJhzpeIt1Kt2qo56K7+pn3kDw9mCXCzaoSOJgjxmAyL6h
Aiy3edF9H3GsbABnN+iJmKLNsHHI2b+pooWPW7rgLGFyqsxA1EU6KPzTayS2n0gDjo0k4qeQxFXj
m+TW8Gk4Qyi5MPOLslLFrVLVKs8lWHg+kmZyvYHUQAklwRfyWEF/HJtmvHZXHEX6nh0ZZhxnHIA1
fS3ChoxV7Fw3nNMzj53V0jU1yh577++C6iQKwfiiJRodPVgnVgyJ8/Hy3spEE8xd/OHC30n6r6J4
Jd0cB5ZDPnyqqvD7eTPzFgUj08+9icLj3Dn3/qrY287Rva2N230Q7KVSLIG3Uc8YEyBVKbslvCV4
M84S1MqEdayA3N3/xuwwc4D0W581FUrzP2rMaZem5VqE2TVoKr3d/SpdyDI7q/5BG7skgmHaOi1e
GeY62kAqECxqjVcOqbCLfeTCogQdkcvpJfL2XhF/7sXcLeEwOqQaFCMAm4CZf5Lb6GphTb6XB4ur
59lwGr5cZwnsSOemSGss7TetMs6k57p82j4rvKU7NfKmHmr5R/HdUWQoJ03VnOCHwa6F0WOjBgAp
L8/4GMvdfM2a0Rc6+e6ke5Y7Hm1oBKqg/km7F5mYhm//LUcMReOd5NEC5VfnIMWFPllAtdjeg771
ZNbU3fcpsAJKHN7jQdaXKnyKyBpxHxhtBUQiNZvCnBi/DMzBCO0f+sk7DMwCjvNvSL3sfKigCtOP
6alIe6Dqko70IjgADXwmRszRNOHfZ7mLJmWIG3Q/veX10TDpzvCF6A8IsWmECByKFtrsDN8Eh39m
6ADPm15w/K2bwi1uwhCk16K1apRl2qbp0YRvH0soEe2FoELWYXIUW1judzGeG62JXw8WXeh0iJDu
R3NgrGfF/z1gcz/vc35i0r4q3lY3tE8UcJvurpVoD2UdVa4UImd8fPD/TFSpLHSaYqiqCPLR3jYu
hqzSPVNRdUIK+9CAAUVPKlpakLDg7VHCKoHjKHRNEM1BIK3C1qwJLNAFLr3kxPiGtTMidfAIM20F
mYByYj2Xm5uN7Jes1u8T0EWpEIjTq5O2lw/y2T43LYbZ4EYGUfLxzFBMwd4bYyHcd/Mp2VxRNREk
bLKXV3o2N9dPXrx754B3D1dr9t7YcuOQ0veXNwqK5LNuAvJQdN/OiCE8Q8EGXMEFq20Q0fzKjGOH
as3BKdXoquwMnurONr0BCjH+dgm+cmez1e4NaWh5QSKSm44bjEo55DAdLo5wjN0VGCs+DwtQtEld
ZPdCetfCfAQuTxlNEMDI3JA9jRITRoqE+WgY6hCklhJ819fe5jOuJpprXM4n8e11PbQWJKOEz/C3
hsCq62z/qjKApZGl9g16ZMW6pXNHR5xnyDHh/CzqRF6aiHq+mTydcScERbr1YjBm6AFJuMawG+Vv
T+cJoPIXHkhe1nEm4cXDoIIbmlUVFYG++IkuRbVuWzdAQRD+bmf6kEwCwXBOlHrDorx73ojsh+ly
T3BR9bglxKRYNBSB6yc8ywzQdhKj/R/EjuHmOsEy72Dv0r06gEvXm0M/kc7dMVUM3v77eGfqkpGz
8nnm8hLW73BrUFM8lbpDrN1b6yH/MmE4j1ykKTeSQraupe8vOiebRppGCXAqeYUl8naC0tfwjIXC
KJldyGnUJq8IByGkir4slKaEz/a3+8/XilifkYxaZWLtwvMktAxC9P6eBQvakxJrizEY5H5djGCu
yJ9mn4IQ1mavSJdnzzbIG1qG2KdOvWsuPg1AqkZ5lSfFUa8MS76EQAaBjToG2+pXgfVkv3Lq7IGg
zhlIaxtHMZp8pjErlFc1sqwiDN8sfNJZ07qNu8m+kfVT4F0oKqbccoLp64V0LQT6c6p8r1+W56dE
C/L4yh4WKOya8JHHc34dVBjtrUtxdEoH0RPtjXiT4R8rbUELr+kVl5mUiEPAIDC6TZIip1BUy6a0
EGpou/mSfH0VXgt1SdGpA46iOP8rgQywVOFrXiCnKUixORaCSSDSjE4PFJ948FidSKIdGnlQoEqA
ZI5islPlEl41y2Lkjnp3h/8OpSCQX6da0qfk4xauBsam+tr1c2/bJFCJGL9YUZpHS7OfhR0i/YNA
LttUbLt/NIkVHHySc2Lg8f2XQUxeBgundCC4FxvdAsCDteTZa4z16W+BPNUe/UA6SGz4V7GNcg8H
8R1at8yfTrRDm1JzmN3ryRBsOKtea/GzhDNU61v0ZKpa0aiv39YUmGk01uI4fi1yGh1qPhHN7rU3
kBbVtRn0PMwbDpA/dvjiOSdfikYrIbWUxPSObYqpYZ2xLyBXAOlAXfCUa+SLFtB2HpOiNreNO+ZB
ciRQuwXjLSizaXYHWrBPjP0at8ABTcAKqlZrhKiFRKNi2O783w/6j2qPeLVUdnnd/+p/8Z15hIQm
d9nyqKGOqV4YMQUaod8wrcsb2C6PslVWUM7ffFKU1wJ8geAUTDjPyVNiotcg5+nlla4DTQqqcW91
wLeyRSCR9N1fbS8W0Pc2/I397eOIdJTOO5tkQvuwzuMoJiBBLDwBm0qeGIbk19G4LTL/5GeVO7ZX
kJlXqeDr7MN0TwKn8tNS8uM+NpjxsZVfgpYY9852rfe+NwB6wy6zh+8o8ydZ5XaVpzvbFVqr+OYI
MsNVpaGvd0EN+sJaAOuMqQPKQ7dtEFc9bakzQZNHajE+mbUYajthWhfreMfZLr48kRGOVsvXVy2P
0GetCRRtbhQIIwieSowY+4wuBrnfQJfj+nLFrXlt9BHE8dbnverJsnjByzhXIji5sINjG/5I7T9N
itwvE4/PqHYK02El25mOTbBmOv1lbQx5a/lTsNb07TsC7nRHk0gm7EN9ExIAKZQTfhicFLQdiVXX
s70jgE8Dgp3Yo8vgjjPAXM71q9jP2z+cqa/ELv+TcxbIU6YLDYtbXt6j2DkDKsaJybhfGbyKm1DS
sSaWo80Umn3Xc8Qe4HFrGO994P6wihwDJPEWxKqjYmd4grAC+7l1b7IOxHx/yu93mhu/ALG0kz32
M0kYVuFTXKNIoxQ759xFrJT5Q7q7ClJ3G2wqCoDNTnsZ39k7zMdgYlakENMcd4tKuOYNEwefL6LV
AjLdyDC8AGJcevmo6ZsnuGJtk39Vn1rnr6BiwSdF97OxAzTR4xr9hz/NIiRSoeqo6gL03keTqVaL
ty6oXdz5kvc2QyYHo4LDpeLYQvOPXBNzF48CujC5x7AQ6lxqEgkJ0Dp/Q4GjgxTa2vF8NtZT815G
/hWSmpKwnuyguhu2MJNpicN8eANyqN5T11ptuZPy4MZ0v/7whHHJiTMOCXGQ77trQAdzmCGrS1zK
kLpsf4d8zg/jszgmev0IU5DBEpPTbMVQZRleg43Hc7iDL2cytnbx9L+cGmkZdCAmu0MZGLytaRRJ
Er3tbDNO8QJFjqlJQPSHT6W9V7JlG0u+RV0UK6nm757QC6hMEQmwwBbiBpJRkQJ9QQBN2mEyGSYI
4SjEIG01j7RsMVbptu7AYv6fGWwyMNQ8zQ0ZS0PnHsh6sGask67YYcwMjtBaQ9N4lOU56uk6HJoI
mcP5xHwzqzn9vQ3+erK6svKW3t65KNzgkTEHjrjIX/gEv55PXSe9VNF+lKJyWtSjp4dSppwujYD8
muSZFlK3pRMl60C6M3Tp5y28bKBrhDpPmPMYjsOBGm46jQvg7jkRAk3nnurYQpu5qC29TY3OOnTY
qvSejTsz/yBxNCrHEPjR7i2k5B7Z5Tgc1iLiErMTu40C1pN1g3nDMTvfv1kVXOjKTtAaUbeZgpgU
p/nJwPX8t4XSyaKUI79zmDiJSm6O5F6p879f8NPiWXUgs/mAlwDas+vxv9HumA2IS7ecN98KD1MJ
f+lGKQRpIhga4PpLthdW8o/EZGEZEs90xa/X5qobgBgTsiRxn8KR/aoY5nut8e+XdcV/gGDUgfZf
22gGADGedPqYEeAgGQqljal4s8bKN8DPLacvRmG2dA3xCpxoDCMTMsdVT2Z2jtD53NQ2/vqIIseN
xrywQw1h5Fc36L/ZQ0Bnh8w4G+bMzfgOvxRvCH/yI0IJ34CioutQBTDxIJ7Pes7ShW+LPI20urSN
g6PbpMhLDxF9Ku1QqhjF9p0BXsJOXrPitKGu2QrmvVN6JYPsZSPoCYoXW3uhROfpJfP59DBlT2DH
JkQKoJUbzeCkIlqg4P69pxQxH5bVx0EJ5l8YBPxppUEc/eHujrV4oO4938Tlq+ZtOE+0LWXnG8VH
LdLLCYxV1cT2RA41Gh8SX+ixgN22jWBz0W/M2j+dqh7lMQc8vrmWRLLayjoQeH4bk9Qcc63nU3we
U9zFArD3twFQ+rfJYjP62tEiYRqBS6d54NwHUiqcIlK0NgXHjIa33WdH6Jnz25xeIQR48KslVmX4
NJpsXKl+qJ9VUrTPJ5p1OkMVX6OxUb3RtoshtgXHdfWzdo9YTQjqAR/jdPEo2WoSEHucPQ84Kk4T
okWitUCAl0/llAF7sGmZwYQu5sejz2Bdw+Bw06/11bcOdNyPMQUKgrZJ6yqNxk+TGGs8BdB4+Vnc
/mCNtTa8FYkubLvznWDNPpFDunse8QPtgaWGX5uT8EWKUngY9YO91YV4hYRIaQK5gwzNxYPjoidm
7YPNGkW+1bpUy7+P+StaJHIvrLllE4N0zAbdyZkyDev8BprmRxHKhaQXjAbF7Gny+NiNRiMU3Jj3
QSXfajJAa/KLRpSV3Q5J9De6rTbvoD6FolG1bpHwFsTJo6PgwbRvBqj6x7pkRfzAUUkSl6CUdSDI
KAwK1tiIpSgWBSYJexHMKYm2L117WmAfigtUcDiY7GEIB/JtAjdKeGN8dlRHe0ZGP13bYORRtock
x0EJmpAEsrttLxsufJjKlmJu/nI8Z0OF0jE1vVTIqdu9Q4Ufgntdriynjage9rc5fneRiwJudztq
5NSBzCZiX6k/EUG/t22bKRUj47W3sPb/68baoRRPac4bt24MoWT2Dm14cHTpOQvATHma5szDog8E
2/syKfY96USwb6oSkIYZzYo7ZKLHHsGWfVOPl32MJck8zBu1uIDU8ScBAlFyc7pOfcy4B3I5/BRe
wAVxsdL1AQAgugPlikkUBOv2x9Iiq6zVaul5fDFVFGE/58DF3uJYv9dNa2huNjnUlCJlNC4kEgGd
kV3q3F5HhIbq8cJucV8NJdw6jol84Hhflku6UmoWkAvU3qp1HxAHPT3nQ5Yd0qJM89a53i8GmTso
j2mXLPYUsA5xuOUjbj97ru7os597NAd1heL1IV5eErTwHo6TATDDEzL/BguvGvkp+lgCm6lzVxsx
Ads+qkWcLI83uX5zX+915F6+MJ8peTKbhepzvQqFSyA7EgXsbQVlPJHtcqW1zRwjiebZUlG9PfWt
gUtdKksnScte+xtfK0yTS3sqFqqOJsDNwS8G1ghr8q5RVzkWv9jgQrU2p1IxvKxP/XBqRUZ7oXTA
rKlUfIYyRm0NqSam+XQznAkl63zvukhBtmXdJku8JP/4UBfjLex6VhIiDteBaPOEKl0MNGkeoohz
OH4BiDu053OcrDxWRBODDCxrOGtYNSF7JrAbtzTE0Z0oIXomoejCYwzAkJy6L0Bw2ZhxrhU5UsYd
rUOKiYuXKJm0gGAzgz6w24X0Z3BKbj5k1X5IwXzrDPlV7z5xhF3dzxSr5rRBY5SHeIKojI8Rh5gb
xNvAZQiRhR4yNAd+yz6Sm2ZtSOHWtsXure0PXkBcP/STKzkmIHecpYZ4nulr41/8YyFhqhm/cadh
xmVu2GNWgPMLzV2tCu1yylUkWIcQD2N+9ycPgA2PsrLdGwwBpkRx721YbEmY8x84Mu64NtIqu/RF
alqg8Lu/xEaWaRYpL3m17qdFs5kytJztObeAWc6YetPHHr8QsKuA0SPlcX1gHFlQtnSDYLP7lND6
/CZ4W9as68TCui/Z14YrhG71vPuzb00jkEwMwqODGS0fAzgin27gdUqFd0zizlZIRgYQGGYMJ8AJ
DNExV//C7u9cE/KkmqB2F/EmSYkeNCrB29XluRWx78oSO256PayISVjhDlSXlr9C00enImA1iUV6
FHt8i+BaVSYJh0UAApFirsDjSo2LXOoTaDcUOw8I+2JX37JseFqDs6eUIC2uTrETEygSeQyYcNBX
dGdJDWDDOPA1/fGFXLAVazRYC0/p2xEgZdX53aQ7mL3E8HhEdkqA/Nskk9IjScNkq05K9uhlhcFm
s5CxmCBZwt23JL7oa/7KXa/DZAqLxOiqubyo9YSk72pwJyD+sePzK0WnwOeSKQPe5MqbCSL2jorw
yw3XK/LkK68DC+aGupUnzmrf8dz3gWZ74nw7M0w5YRTqIpOzTCZlOnmuv1OfZX8DueCMD+M36Pd4
r0HW8GgjZCSgs5AEaspHGn7KCFkE0W2T042ZdiinqngXt1PVPjzmLNBVo21P+9PJ09RTsecakKBh
M8Ih8GAT6DlnnnM6XWfAmC2QcJzEh0bx5Q2HG34yLDvuCG0MoWevAm2Y3qKhLv88PZmgQ0A0/ZJV
JKOxMIFRIX5fzaYu6LDoMCDjsXzdJtFThVR2sGRPWswLkq9aEAvWzml5vmTXDZb3+xLey9GqPExw
piYctFGs8ch1RVSnUNrPmmrMvzEwwGXwR+5+ZR06SdML0gyt0S3EVm51jvY37J29iFWgcUSPl+Lp
Bdf9JKA6g1hTV8iAe3jMx/VIJzMJb6EHVscAHI2TPFVCFpOz22v0v29At9Cdl43dBWWiNPan0r1t
714u9fP2bwhdMBftBja0tzFp2k/p17hWWTKWcSc7fUVLg/KqzhJXl78eznSlcZR/qFU7iqt/p1FR
9bOQpZCeBHXKXCnQDnDtuXW+6ruVQXOF1+dv+lAK+uwHiD6xcnL7boYW9PWRULuM7LiyuHmjTlfO
WSxub+5mkkDOB7y/no0ln+akmjt1w7gZFyMPatCFoqV/T7FcRekUkPnxKZuGAwyekSqqMd1GLAVZ
fw1FlDB8FKPOUt135NnwK664dfVeYfQKYDu33AXZoxx242/7u4Nn3mVQKgtVIzYvI0gsey0cZSP8
oGHwyKOyJceOyDgFjvp4eaCKhveyDxMV1gYoKLxs1uF2zVc7ET3CjxPzYzu698noYT43uY2g0pLW
q374jpSNFQ5/l9iPEeZkuZ2N6sd+2yS+EBeyDNScPmUUZLRoJXdStsRDl3grhiMZADx1EeBwAhnh
MyupUTo7xoVqaU7F4j7zaazzbSdodMGWAIipHKMLnqrhjyYeOiAYoAOmmNauNvnGw46GH13hIiOO
oP43PlKYJf6dSwkd+iIxNk6bOgXl6zfXMzAYoyiKRYASjGTS/cwCF9GTF/LzZDrTzlvgkU67LC2J
OvWLVrRDm/NYGWplKjVYzYUkd3JA7eXJ6ufVIjTy6y0XJNK5/eE8UWMi8SSaJZOGxvDQJdaerfnB
hy+D3V0fwjV/r10Ao1QxrslE9BqwqMDQtSRtM3rFMxUqI/BzzjZrbOppO/acKq55RCYuQuKDkGQ7
R0Mpce2SaIN2zbskhD/+NpGsbskIe+zLnxbmVXPQzw8xEQLNcDSaxzDF+bxOeDn2nnHxZTGoGsbw
AYaqrm3rc5CJyZeyBn7txzcAhMraLh20wg5SvzvAg7tS79IjL3uescjC9iJr/rgwAjyeYfW3baHj
6PcZYwSjG4zv/NHyrCzeFKlF9aPu9BK2Nqsn4fhwY+pB0G/84XKldTDXZvGqi6h9NsQ+1x0cs6Xd
SUiRgQIfFxl+y/qhI41DEyqtit4y9a45s1QykH1J2WcGDfKXY/IjWjaPv33DZAfNEl0tzpu07XYd
eyV+emzGrlrhZJxqbSxg5WPC5//iVGgPMRhXRfwaig+pdgo2Mz3WoCN9pKGH0u8gJx9zXB6v/ssb
1wIqQXOzMILn8hD5rtS5PiZp0Dy3O7xVlfQCkbQdunat/5TNUvhydMlpbxkiuetxLxQQUeW6BfOK
NzHGOWzX+QPGtPlpy7lwr3gotLAMP2PmX5HjkxSRGAWxh7JvagbZKWz8Jmcj1p8f1S/7P2TB/wvR
/m5V9T+fGzqKPYaygmD2x8TkC0ZkaEzM6Vi45RrGWUWOMd7d+F8MfF5K1+r6F0lVevwwhZlrt7Ql
Z75u69LRBboV4bbQwlMhXlRIhd4Z5TJ9FXdNalGUqzPuYoxsqdSkFFTZfGcGUzudCRjnSseydAsj
wUQycvaK/6yHu27gfvhztqEuYijO1cDCvrbx20EnipVu3pP16Hy/Zi1jNQOocR8ieKIHzpfJejES
8UFaYsgbvtKoWvcUTIk6Z6ENtKjtZZm1VSFdjkSf611Wzv8ivETS+O4shn++j781BCp9KOBYlkTR
MWGbcm53+cPMzve3qN72pcxCZibDUWU46cz5c46V3v0d4CPbD8bd6hXTUj2xRJ92tH84LIG1lrB2
Igep7RMOJEtXDjQA8KbteL+pBLbtZ6QadRcVwQYIX6Z6u3wEhWizLrMzE4+zYUejpclALkx9irrz
+F5572i1yzNQgpC4+Zy1pUYWsS7Tqleb7dbSBxitsRaI8JksGUMOdlooXehu2k050uHmEzqQ/cHG
YlKRYafOy7ZMXEeGnkIokjCEnkWyO4288vB6C/s0etwhjEtH6h58nGoREj72qXOPlZBqKGHHgiPx
2Ov74vNkpwxx080ZPjmEdOwCXIdu6LEIJVclDfkHCwwuI564ctghKIzvo14s6VUrx/0Q7pIiOZ67
+q3t21lSDHfcWjmcvjW2Cs9StgqSRE50nqtB854w0Yxi+RCm0+FAPk/Y0kiFo99RURQUQwI8vS1+
pIda66kJ+1FCFR2RCsA9hoDXfoptv3tW24M8FekXEBSe1O/DRQfEqcUt0RBMYB+sznq30pkJK8S5
xgzfymVuow/erBO/YZb1SF6I9KGrwy14WzobmQjpU3fca0w8qWZcmx2n3ywJsyyf/wbXwwXFHe95
HT0pp1OrGqMtrXb/nGZSZyZjbTc8eCgQYkq+3HyQ9thxjUhsFoZyRecUWe3o0ss8lwGPQzKIr0xi
46jy8A/WTYWE0eROjN6IrjosGtTnlSF9h2PcRMO+2vqFXsHPCvViiPVN5qxYKz/KL3joP1Dn3DDN
UobaaYmtC+6dQgRpcNBMKCmdLWstZtKWIE+6DWZNMxjd9cbZXpj+Syz6pDLg4l5BRu/WfweSVotA
TEazpEWgbLGmO1zSQ6gmAU3XuDR/L9GKVAg3jfskRjPMISoTZhUnD344mkx9FxpWuTxpPjomEQR8
jy5nrejPj1FD4+yTxX6NeoO5eVCOqZuYFfQbS3A6YXC8uLaw5kwrNsxB7s5zOmfz4TqGn1zl81rv
rtJ2K2dBZA/6086SwSJuXhHbuyYMZFaUO4faYZnMR9R654dnwb6B4Jr3YiRqN0XggXYPG9kCwL4w
Tgweb/p/YGNrSQSNZFHNejle2M8J05MhSrzj/5t1cFDqD6CaESVqTi82Lc3cY74LWWSQxkL+l2HG
8SeZkzfNPL6yY18yQFSQpLK4J41Rk+9fOUtf1F5eFMvYNN5Sx9Xlh70f7bKU02RTdUUTxLKZTBIM
aEmEUQwYMVfv8FAYOjsBsxUU7xv3c9sD0lYbl+eOr6yBUvR0/AuOTV637Dx4y5OIs0iHyZKbYZeD
8RetnlpAJPSRKCoAwxeghDES3kj7pdfArFyLEec3ZItvT8cKpHIhhW6VXJWIaZeFnN0lEiHsVBfy
4I+Gb4niVUK3qpArLgm2b+K1hPo2JUlXZw8oSiwIURabXAGWRvOfxWNOpabEQniLik5rsrCTaKGj
ZXfBRHwYzkglhXSjL/pHL0Me60AD9TzVgNPOeQYvHn2v0y+5osQSHScle3OBItVNie2f9hGLsTNl
WKxlcYzNH8oOtOXsKiD/R+0vGml4mrQGSWYElB2hc8DEdrt98dBSgHJqYv9UT8cKzuTgl+wzAK9G
QaD+gQUqpNsYontU0VV9fqfXiWSdRVMUXTd1N9fZeTgXZcGcld4+3O6z5uHPJrGujGkvEVOPLVth
/GSSTjry2uPtcUoZKHKiNx2EEI6GK0gth0FD/ft+bxTWMeyfAtK6xxN2TcLyZ9CCDbHTVk7cEgvj
s/JfWbrV18f5UlCGsE+s6k1xdaP7D+3qYZst7dzedVcBVU3pvAwWTHWSvb2Y6oPKMWEcSVb5YRq4
QbpjrClOdLa2lwFdj484BmL99n2a35tOB4UKzA6b3Fsjdh0F/To/PjaOw2qv6kV9OGV8o6LLQdVw
3CWMwQUTopA+Fn93rmXrd9YMFxP9vELelqE3FP5dp2XZ2Vlf5etJQ3iLt1WIoF9UuqBA58+EgE9J
cM3LQRYIkxhRDjzwd0b+5wmTHROXBi9HS3FY4HpNPsBo4rUISD6p5tQB9bTJ9ju+oagk2lAencJN
H2mDgof2xEST/CWAo/fP9PwToRi9wQoO71FubRTD33UnAzCgvCEj7RwAtSwwma0g4XVx/p/BSMLd
gp7Yj9XlaJVXflN3dqgctHqnlS+0F9Jd633L3SU6Sb+/vZayOxu2VlLnxLvcTHOtbzc3XUMM4z86
7R3bYRJHrwkyUlTAtwTGR3kEEJBsZCK+E3aV8U8xFIGvX249HhcALAum8Uf/cjKzuI7OBdlg488q
304N3FWMfKV9JfhNB0DaTQpOHdpSqfddQy0mg7MQ/bMhjvBMfdKnmNlKwZGLrkSWgR3JyXCFeOrl
xmeUy+81yT2TOlSbQnmo5IMCVnQW9RlXK8sUw9CLDAI5PfZVawgJh58QoDIblEbGu+MOT4S1JhO0
VeQlrzYHP1KNP58oX65E0gW9Uubp6Y+VTykNqwZseBH7HMGVPilfmkXfo7wQ65AsSPyAxP9SIWYE
kEK62AHcLI8XSHrPSvVO6G4Q5PWDkVfiC/PJbeSYvVTo9YB3PB8Bh28ji69i4vsBS7PM1CHx4OlP
IShrVAnaWLNnk08dbKvjilvjlOv96JDRznXDqAKM4gnLtQf4zmt6vdVaEBYY50V8nCI9heGjJlcG
foEqvl0JLWh8rKkxSsRVek9NNOfDOeuP35aYMsUaJiUhRWPyGvciGusOfOK0EwyU6DvWsxGhvd6v
xvKWsjD/Q85NEheFf8wCI1c6hzTwls5K8d2ld8N7LXhYV7wbqOG2cwf3kmN99EVfOG4pjXuhk40j
NWqY5+eW94spiPeOHsRQokOe+snCnpJZTVhX3FIfd8KlgmOTE6TunQbERRprFuoyZrVqcYsUZByr
4JcCHExdMgCyvRnrcmh3LKBdvq8Ajnxi3mc1LM+fKxPKruSCDptuDBgimI0wbraTeYyf9f7wQekg
Y0uef3iWAlldERBbYzISy2s3iZ7SA6r4hL5R0KKwr/kIsQrjnwoiH5AAAQdBMgQReANsR/gRRBCH
tKiqeeUcIz5ukqo9aSFi7+tLwv0w3GkrdZzYAIlxYjWKHLjMxPoi6ED0MXIOq1tUNyAP7wf4G5QC
1F9bnz2CWxnsHbSF03QpglDOrR04lWiodS4DSw8aU5cTVqi3s6xmuZuUAgeBKJ+LHuLadpf9F/kX
YZ70iL7U7g0RZuzW8MmJCOVuZzvMZPFaOl6nIZJfGi3CwZsWrvN642SMxBpH5UUq9oPddAYJSL4F
c/GbNizH6lSxdI00kiHFFGumrhJ1N1bTsv2GTvOI2S2ti9FiYMHAj5pHTHUt3B68FMyz1zyiPuGd
G3NUFAP0/CgJz4XV+ZnxtF7BzTFqJobvYrpx+qMx3xrTlaqdn0hhwQgEJW2xxZi1SgjJ5u/mvqF2
3CXMP1qUycjUsRpeTcimR40g1bLqZ6CJS3lNqAhZU2I7btzty+NJAkDmRv77zvnovUSs98upzFW7
RfX+N1nOBF+vIr5su3upxaDASJ1wsicul4zu/BwINv3WawWVdt2NzZ1AX2ngQJtCvxwbEpIXBTW8
UKQ5fTvLhljb70NHZ1rU6EdYKkltbgdpnQ6WEjW1E0TfmU0feKHZ6a3YY00gGN84WKmhPjg+n7Me
C+pVB0ey+06pFKEIV7oNI5OpLpSiEsE30iTG4kx4Tj/OXosJjpRh5f0F2EgesrLcGad2ET6CgiEk
t4R8Un3CoRVX/9k3eDTx8bieMrOkQIzvPW9FI+DvAucAZVCjsrkYoNUTeEZWEk92SrWiBdkmnuni
g6S1NrPu+9sS6jduLyQOuS6hwvkixuGHKTE9rugwPhZeGqaaQ32Q9wlZ+Flqq3vvh6DmcGXw+JYf
MZkKcMY+O3Q9ifyWOe5qPb9meAdFxNkSNed46WFrnHBsvjBA9MD+tonXuW52wOTLvtnW59PUYxRq
p0SNEcyK222bYEJR1M7mlqi816bHFx3iUBoCGKOtL6ea2TkozdFGBIiODzy+Ci9fK2kIcSS0wvuU
CysS69hOybaJnoRAgojmpT9YVkbYaDK1gmq6eEc3121Azu7of3ksFgvB2FVXPB4mz7xJh9djaxfV
6FQwq38Y3IV2cUK31d1Yb21t+ZPnsYoOH8OINcmvEmDH3Px9UcH2kbxweLA95hT78o69/Mo0ukUm
zU42OSg3hJUjwz40y53eI5GXdYSq9oy8VA5SRsA0aRW6ecm4S8DNw0BSRyTaDsvgrbAwAFUw1/5P
VHxeiID573g/CNsS7doNBc88oHid1oQP6yGe9boDdmq07PZCl2agybhuAWmpW8MCR4XGg9gYyuYO
6fdT03P7Cd2dCXKuSzNOIhoz1ohd3qsDqUYy3ZoyzqvpbxV6/GIvNech/fq//CXnlbreG0ZkN3gd
IPn6avYL4cm+3Pbc+k2vcYh7bHtvKQ7CbuV+6eCHC3n19NwF9daNTGDiuHsUdxfpXujabuioDEUu
+WrjYRuljwGqhcPcwhOwMLvJ8+dR0Z0Prhk/Zzc8ZUHpWzj2YDPTvNYR6uguuzs3cGZTlxwUBDrE
GaY73yNDp4ClsJR1MtSykFulk88kz8Rmh8ZKX+0dyizb0iHGlkCDoUKGLqwnLrMZ70a1gDdBrFZ5
dbymI4I+0CqwL1+CwEoSYTFg/NqvBbE5rUlLV2EyRdhfM2hvvwpuz5OvvlxhizwkWwHdBt6umxPZ
Io3TBr1tkigInaNHb6ZUB2TQE6sDRREnaOghYnlDaqHUTj0QSpM6ws9PXcyWZDrnTbbMJMW9XPPZ
nMX5obDs3hLqrejVnsXLMgJgz5r5iyPRjz7U/NOqc4J5ubGHK7Ukr0UXmxgkhGndrBIsAFjS9vGN
5/YkT357gF0rMHulD9WcPQ/4JUrABO5F7Xjwe0BmlUAF/N48YgCIYCRGLIH44gvoteSp3NjtFwhh
FtFuddo4IajaQI/6KYeY4ZRG8xqPgByvtPXRH/OZNvV7iaeRE0x4XDNEfGz0Dq9tp1lmIyZj32cs
l5y7jHyNpx5w+zor0MMAtK1SJ5189gIb/hGeZeI6niZ4WprdxbN2UukHoOV7ux6nelmFhRG40kDd
g9+r2f92WXrIFLqcPyRQoVynEWhzVwT0CwRUXRJpeIYdSQsdseT/4gleSlnMPvEu58PTbxbq2ism
HUToRLpJoF7kj52EtR+OCvkEwjZoJvh81ponPbYy+YHp03NZJO9l0+fFxslrM6vpJuLXaMXc0zVy
K8cIc8mPQsERHoQDVSxScEYKpZrRpBEiRPs32pJbIgFAEaBNmFKo+m2Pz/7Wnup8ua+azCRghKZu
q8Fo2XqVWrV5nIChWaJtDXo+Id8uqzFvPO+iF/5GN6g6ypnWzlxzmRSf8Wcu1ycPFLtYlsWlp0+a
z7MmrK+APUxyRVDa4J33pDR8topa8n0wCOHE4SCCyZjLFOU00yDC9kwhzL6B2or0Q6tDnF2V8Hdd
uxmTBdSkH6Dau75VrpWjKiH8ZWW9nkbgOAdolQA3IU2905jlRPuTW0wCOuRwWvjT9iRtWOsupT/+
vPk+Zc4/Xw8mQKldc92q4i7b3eK691pCAHEyntzVqwJY6c3PmU6W/H1x/2RKtCVrFfa+R10SxNPS
bkxTjZeH6Qtq9Y2edDA+aprAd2OsHd5+grwnK61IgBL4VVot6w9LXKesa6GtWI6aJG3DmJeEgJRb
dYj5rmvZka2PgBBar+qye6cBWzDc1oYDkk4zOGA+9GOW+QrPLbLjzRfjrOgqI5uPqw0zD8v8Qfc2
ICefc5sjHiH3EVxA9SdunseY6dKgBn0CPhN17gu/GidzzreXbVP8qzQ62w5gve77yc0+37ZUoP60
0AwBkx08/7y0Ppm6cYVJu9BZuTV068/RHIWNj1Jt/yokS+e7VjiEpHPPqtmn0BO+NHTyrAzkAh7C
TJEiImpc5z1lQqVri4gG3TUF6xqNB8dBwQUV3ZhHKGw89ZzVfQ/ZH0s6xQIXRSy1QYzrCUUGOCJ6
VsiORBog493H2LSmNvAB/yMP1GhWAQeGyrFEfFariagNQthlWayfOm2+A/CMgCG6hTl75h8gg/UQ
+a3vAe+3szMnu5RjD17pTsAXqkXpZ5L267jB8kwyuQDq+b+yut9/yisjPjni/Zbk3kd4ORUHX+zl
woQoUNy0JHnPzL++b2mxbxfS0wAwbfs/srX2OM/5xIg9o8t17Pb5jjZGk5vuli4Kle4r5U+dCERM
4u8N12uRSArPmAg2beqHniiAxUlkiEa3GOi8mRp6OXHu+PB/pd2MXvgVaM5mwq6+5xKAEfxa79OB
CethZmM49DgrlmTgEEqioM7W4sFA4wIL839QyYUHsiizurjPXk6tRqlDxfHRSuY6U6QAzZIvlo9W
P6rIZCDpQ9ezAFiJnNLTiJQRJ8lsuZIVOmtah3VZuXoIj/5z3AQpHslvWV9UDzGnK2S+9f7bN1wg
M7JJtt7EtsooPIhPDOnqPeZMx9uoELSoXY2HHxxYIddNjf2koN+jkeV0u3CnztLj9I2BKPrAzro3
yRkMK9ehPohV/TE38wyN0Ii7ry0p9Ah8UcQBPYwmWxZ3ftO0RIOZ5jIiZRYqkyM8QjkeURSvvfNa
QOcw6NYdwHH6dt5/biButkEC6VQ9XdfR7IFnyK9aKfE7VnB+5FMnIuhKAeeFLRvJSqeoc5a6+xv5
ECWeX2Lh0FiqT9yEbreBc6G5ESYzql4KAG/wL5D6nsmayOg9c8Wh2RtjFI25j8dkTbBQfUIHFy2o
nZdbTvIFhG/Z6nPqz/OAEGjIEmwWm3TaixFmUPVki5F2woCohan64x+ddxUryWDV9Y+biecluVCD
a0foOttocQxPmtL9sYsW8gsJhNPBGCwoqQ9vPWdJ38R8p1p7zuPhPt1JQt4C8739Q+7zRh5vFMhm
m2w66wM6xNDcV3fSyKjO4pLDm9PKNNdRn9RaMUFNcqMuCZxmLcivpHSf+8/SBn8QwbnrzU3TJbu6
8oxVvnO4Y6CuAY5Mg7X00quk50vVGbO4iQFgSOgpAYUWbaL5FQSrITjib20j6kmI+CVXIBxdCawy
HqWwd4IGemqNuPMWEIC08DIrgrJxzt6bOMEz9zcpQNUcrzH6b7U7L7u7Pvf3YrPcACqBGOOJF41E
OoqEnb4PU8HgpP2oSZFMVIZ+ItjAERGQRV1xQFo9NVHdBhbt4NkD7LHe09PhLcXOL06foZpEK6S4
s3lQF1TvOnCWkC4Ujxo68a6y62Wkbuw+lKsGy8t/uHsRSMKXViPLS2PieDPZS3yhuGRXkce9hDTY
TVudlvY8gu/49TCI4vqRdRp0BO+Qu6RtABcEAMAytDsQ2Iw0FnqOW80wFAZHQYJVUCCB1AzyBcHE
gvKTVEQqLcJJBgkJA7hNf+s4gpxRi8mYCf9+1yBsbZQ++wRurFxc7+skInxVkzYRsNoOnKXP1wix
odRjwCR+BIOLY4YUWxohtQsYZSNfZ75OEzT+QTBog6gB+ayCunBeu7w5PKOGsntWyAZtm2Xge5w0
sPX0eKp/A8AzNxc7LzCivduA4pGJL55NQ5hEnf3M/MLbeO5hqBACMtIlPniwK6GuY10B8X5NrxvZ
wqHzR+qkdJRdT5k91Nb4bINT/559GvIFd5xclg/wgFzHi1LZpepTiW1gdKnvt7cY1q9Njkux4N+H
hMHL4I96cWU3+YL9RXYInaf/jQKoOZGChlvcXu2VWesSj2IJPwE+0DQ0YpM5xGHyEZLq9X+hlmPk
EaWIN7JiMkLcY6jRsKckOuGtwfm6NGqN/CJh6EgxFRtW/6aVFXrvQMOpD5yY6Uuf1aK1voFX2fdr
wl7CkVLesqiPHhoGpeNdsM2YYNQXuQUn
`protect end_protected
