`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SSoBChMKSFCsFOtYbmJr6u9lmp017vqwNBg2ZvVmqj15uYSOcs83IyC0Oz4u8pQhUm82kji4ddZp
/KSpWoFB5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dDaNY/QSilEIHouTSXV5fecvca+JgcQPOGnUWxgZ8Lgzt5nEhWYUmcI4IuVr15gY/T7wPecfQgEn
ZPnTOgHb/pDoGiJj4ordhxgrJrGPg9MkMzCb537uzdqCBFGToubclsfyuSkKKuD3q7XEKszPuCQI
cQuq8rw5hTpNdWxZM10=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3l4BVLePOSQs1rhbTlq7MjbARE/6Mc15niiy1nxu1J/FXxXiaRWxHiLigyt1YuCwj5fn2oXjEVMc
kdzKDhkBAtN6O9CSzN9Jn68IOSsF566JHGbsG8PW5YS88Lgd/dijIs4Bm4FciRx32XkCk8NYShsr
/xOfmXYfmTFYyfz6ziU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rrHZmd6w/oI+5G46Z8BcQ4qUgN7fhriHm5niCP7Vbegd/xYrOUf2kdzcFAUzfvVybsmsrjAvn8aF
z0yMA0LUdg9Swy3gbZ9nu4qX5zXHyJn9+NsZj+o5Wdit5p7paXgGfYQJWh4qI8FMPXlUKb2KUPLZ
P11aEAT9l3e1I9faiJM3UP5uIndnrLhofpoiyEi0anE0IiDICODr4o4NTa9MKOSV4Snp7Zr80wKn
19e17ZxJ3HKbdExWT5X6aBBZq53weIRweRGLPrb9G0Rm+mcek2SGcf2gqVgNafh9pLhKXLBfkyis
AJ7kSNMEQQUHmXaapDR1hcpxPEfOfA0iOKdGgw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FIMJyZfbRqYCCvJI/ADSqIO5yJfRGPJ+hQYeG2Xqs/qEd/BdR9T4AN4a3sT/ogOqCBMV38F0E8b+
Tg09QFycd4dX15etPJgBxCQP5c3cu7ys1UOkrXRfAKXV/jquyLemyVwS2wAjDFV40gQ/YSFQb42v
eKRMqXPVnU/vPgjxuVSrVUm5P/NYSXJJbIlrYci1Vzwipdq2Teb60ORACtG6nux/QfJdP+ASdAbv
3cTvdNbKGykWvEzGAtQNDXKdEpw9blJLARg4pj8kzv9C8XM6ksfTDWVe0fi3TgN+oRsnkh0vAMDi
Sf+H14XFN8/fa6gPLwaZ5NmQGSqOazi/Uh+1pg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I6OjQ+j7PE/9HOjGKGaUPH2tlI4jFYdUAqEwrYmnefZlkXYOCl34I7kwTYEUehz3G+02bUIowfWD
fbUpKkWVr2fwRvTA/Rh5Hr/VFvFXtPZ9G9bRFBfU8Aflc47VjKsA1WDu6mgSLpc8k1E6ptm1g3Xj
LzkGfUCMMXRfP3HW/X3r7ampixTlkbCooODmqzIpSPbxvh0bGZttT2XSvJ7igW5M51c+Jcpog67F
fV95RfXVDE4rWS3bhBi8ocA4uul3FvoJrAa75bRwOATpr35NhPNpn9d7ejhK8mlrnk4r2/7aonp0
CIarND9Wishl+tk1UC1BcWKDsDQYkkZjv2Zh1A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261312)
`protect data_block
HRf1MxbM3/PhIOUHkYVyXkLGDA+4YoFhozHCml/GvKoXEwjJ/ZgXHkWUYnR7zq8EFbHB0m32RyDO
xBrfrJMdcSjPGKdxsNGscmxFFsVf3ClQPCGhlPzQb3B3Qogdsq95y9Wj1LXTXrGkJPAis9TPa3SW
eeVZWzWaMM+IyzuNHYHFzs+wXavU80NRgmJ6CoE4Aqnz1yaXjpg8hQhVhCtPYtvWQTOG/EU9zN/P
XwvtnyAFwMBLbe/RHx59Bqtpz3VxcTD2DdqlLnku3lrpkMAMM/RNALfgUgc4IeJyK442vWzl22g8
k/AhF6DoHXTLgQS64nb6YJQkqZjN1VAcr5Z5nbamfFayXAQKHOh0OYr0uQyPogz/HDAAFHQuUWUW
UBe+6eaChL/N8/Vu1vp3nnM+3huheDF9J9Us1zWHaIPJkfzvNIO0oY5Nlk6mpGKf1VtvDmmnkyLD
YF1MhgM10vUd5z0/oLtAzHqI4xS25BVuWa/PvkUiNNbqofJoPr5KaX1ggAq+ImevJFVHAwO1Bydt
YyNWQWzEj4FGv01azzxO/I6FCAKAb3CUcHgptSFsRw2YR9PRcRwCjzqS0+SigkLzU8xzzfl8h3RS
4rNT8tU/WOPSTk+MEC67BHiD89JVKxi/2+yIQzDvex5duSoJePNrJDGbemaW6TYmcHmO45jhNyv7
vMv78t+tmt5ofs4ImLiCBXTComb1TNPLnWFnL9ady0YEUG2cPeY7hn8V9QWmLtUgqPN4vZ+1LAyE
aNL770ZdSrNF7UtKL5n5OhU99CWdUgQSKfOFg4eqx9BuEfBXJ0l31iU+YtZq6aIqTqRBvVm0giPy
Wf/TvqbZloewHzgtH1m9DY1+zYvKGrXpPAzHHEsg1c5NcQd1y48IufgHjIjxChcqGh1nV8bqREr9
fiJOA+LINfbO6fEuKQEF4Vpys2nGwLvfcG4BIwdZTU1meRGbf2vjdgivsJBDaHJXm/3Rn7lHvMH0
9kyQQcDDkdxpicQ5VTDFTac0mnQsSmNxPNrm9z5g4JWMI1xe9z1qdr3FBLfNULpSdQ9rMuDVDfBJ
PjvKbzdTgG4N+Hp6Yr3B3hijfbqWLELZ8TkotExgyceTK7u8wLvBUHKTy9asYC2MpJuoj0WD3vzA
RRKykobV5ui4HMVM6zZ3eSABMHiKpYwQ9dX2pefY6ObJKHSy/UyDo8YqGSuk9OnQfXxXgowHF88D
0mC6MKFG8vwdFhlSr2p6KjZOAWYc1ubxQ4AfYRbDwODxq0XNZJ9NrA/SB7iO3EOyXfTIBPqhrsgn
C/ERrjL4j9X0PzJ1tmZ0KzTLDGg7VODqrUw+vd8mq22gJLNpcr+AHmGWABXvpuD+U66jTCbjSOyT
kgkc8yO11VZ4FO/9MMyhyKEcca68FoiTzp2L0mCFJpZ0/O1RYSYWTCCmgLA4L2fgI6ous/rO0+Vb
6a1rV6rcLC99HgigWYbKZxZNfgvHQlLnl5eJpkwh4NysDyyanZzpQ3JW0tEqKMmUzQzJRWhNbzgt
RSL8QCcYvajLy9tjS3x01J73cz7VlpMer8ffwbK+zdadOcAVzD9eOZKpryl9RSDwJmCaecYGTX7r
/Vj7Q4KxUMDBINNmwyEXKoqqnx5STvKwkogDLEq0qJD1VpU6bsLqiUedRUeoPts9E2MwCQIriMuj
rU8e/Gh53On+saqD0zvOZ4UulgoUUFgykQs5VMItW581M8TzA2/UkjwZAKR9mLOAu4SZD11acUPd
5FSDrKN5dyJlh+1YpZ0dQKNQBAVIFXFjM3WVHLuXdftbzJJyFRgCldPdanUjAIVOV5L3yK6CmD1f
jAIrqW9BI4YV1fJgOyawad5rMjlDurxObwMwve3R/hbrok6n587q4tobuX50MPVDwSPc2eRu8X98
0W9SZ3vaz4bqmQeG/9u3u5/3pw+Hme/JUYvjYVfkOiAwmQ6CUjS84IPE6/IXnzk6YbFbBcIIaynY
OOCU3xzgG3UF6SNTGsrxwR/G8bWo5krJ/y4/M7POt0aqODGODnVJh7eM4tz3jgoSOlJpi1Ppxj/f
/015rM3ZW2OUriKvORm3Us1ePmTJj1K7CXTSayZyf5HiIUBEvtPMntHdPRBoZDnkkJpmbs0GHwTR
A+iysoRdomKOIC5WnaNz6NKngO8eCzcIm2eO71t+miT3/doUi/TBduHcJYJXFkU2IvRRMrSN51WC
e0tdGAbAGqOkEIBTIW40ZFAsnWDfsJkL1FIGWWrqv+8N8MArSy9E+xxIWu8TL0G70mVuKHl6/kOT
nagR2+J+51uXfpR//JHhyhBRehoRQdac9CwowGD8MLLHx0hAwcVqlBjoVESEASuQrYjS8txSqaU4
iWv+VBeCYyMX3+iMRvjDq6Dkh+nUsTDhpwpKIFPqZ/ba/2VUPfbIkAug4bvpYCPlIGQyWFeW2HWA
I52ABJJymxPhSmMkvQPNexIJJuaenSkjj4oYdvQTuVdQDX2ppvc0+PMiGTpnSrQEFeLccfIWWXOI
SIz6rnZW2vDaZrR0i69h+wuvSmEM4MvC7K5BtdoRplCuEB9B2gSswVY7dFXjG0wxaZ186mojnuhn
ERiTWfu2hyF1hlbMOO6h4/cIYtdhlOvma26YLrUMe3iTUbJVSZdmPRek83rCQKy8JoSTGNOcBHAv
ELkUqfNWG4HIl7rdQWHX+yRUTDJdPvdvmzX2hmMi00krHxKSlRCbExeuKjOn/GU+J81Vxrw02xJO
hty+1a2GXW/4DQ5PcXsBLhgeCrFDJdSk+1OK7FZOwUvcawpKtYOEGi9os2zVIz40zbz21XRLf1gJ
Sa3AyCC2RpA15eJ0XFPx2caGwGBt4KlCyZdw9Na6e9Q5UvzfWrqHlzhdY3kiBhrkjH50eEzAFmIt
VDSyWfpsmbJ06aS8lLW2lRPTcx0dKeju+jJZG7CzDayvUS7gJmX0+dGJXVhF+aJBYz9IIw2vFkmm
sHXMmybwnGdS+QPFKA+U0Kosw4hJ90fbqxAh7+IEo+gYMUQ5tMx34wnhvyEieWmH4zoXYwJpfCVE
IuQ167ZjqVO1xIja62D2G1Wk/LkdRYt60SY3REfDqvdWALm9CcEl5PjHFtdIS40YxzcNt5q2AEx4
lWJduQuOd4QcI4ewiDiNOECRbRElBsCDriGTdueKQlN1KdDjJ4cjynIwAVYHNqOUZSW/nbOS7Qc2
GaAQHf9YrJR6tLovv0CrCZWKuA09/hN27v62GOfqWGb4HUhoKP7vORgNBKcksALYXEqbJI7d3TH0
ijXs+uqiC81T473PDzdf//ow6ly/2uy8xaM0uhRPdWAKE5ap2B01AmtoLb2Q93qqETf/jApF17ER
O4++2Sqli933a9Sw/QQJRFQJDTlz1+BI5lwE8UsirnHjydEKWwDXqwOso2vcY8FjZEVw/CNfyq5W
+RA4g8R3KFU5rCQ8LT505f1/6OwF1qaYLfAtuc88TDcPSGVxesCMA9/jpfRpm08Qauc8BMJ1PhRs
dn0s0SLmR5A7tgTco5FtmQZQWKBfr9G5ERi2gBUlrn/ehSQIWmpt3NnqLshZSBXNkMij0Y4nnFGh
SSTZUfc52y1+fIIW5/0G4+06MbA0bTcT7QB2+YwbTBhLb8vpWv7EYpaLkU71uDiGTkuKfegJVPfS
G1Wjtiw+gbpsD6Bnoysc6KoOJ0RVytU00GLFtQFe/I1/FhcBHKYZEHwWw5YCsnIogJyaev29i930
4nT2tXD29khkZut2RbjXC7xdeXYjK6nPSgQ06Ujjfe0QQ/ZSwC8eLOSP9tDZrrOHjcV4QhmLBC7j
FxSawI9HIC8YoKy5/4itl8S8YTSjbivmuoD+H10NNxRtPCYL4Pl5PxT1ASVHsauzfVAJ+WpDobCa
s12hZ7YAiS2klCpZMyuLzoHcjQ+BTrqLpBuUpilAcx2SqXohTjnBhQjBCrloG4bJTDXnnukEMXjr
z3ZJJnW2XZH3zlpQKiXhPYpKJ1Odtdgg51/GR8c+8SvHHXJwiqmrGmcwue/8WwgDyNA5Am2hYZ8x
oWz8brv+I/fMD1tKJoiJI02RNXJUmvhytNgK91wLwnUNPKFmInrnJmY77essjhQkhFDeC8ITxjRW
RYnTUPisGxkGni4RXCUbPu2tCsaM89CBC3SYslWAZg4sUkO80jYcXMJfNzOVOMbJD+dcCjFzy9dW
WLmw38qb+wy5gUQJ0RpNOWWpoTkarpOK66WstLUVpEH+CmNIPQoh5aiK7VyWOQ5SVUvmbeHTUoWY
hj/dI0U9j/gODOwyQd3k3SRRXJqaY6qVQQtqUutsb+I9nupeew/gZmsLdpHJKjddMdT1GK9MSnba
q2jQSExEMnvBP0sDqo/nXZ4e6VvCALU+FVO+x1dBSDCO4YtRQQ8odPzdQEKPHFTG1SLT+QONJdTt
MWzHdolRF5+HVFuVHC4tjVGjMyNKSh2rT/we2YsjI5s0wr1xa2BdA11T/xNcLvi+myTdyOofAC9h
3mxBwYk3+v+HSRKF1EsaSPB+ktg9j/6yyFrgVWQyhvIMTCLINtwD6K759UAG5kfha7U5JjmlwMU9
YMD8cz4Z1cucQHOQt4AjLHAJcQfxGtdRhvuxK8rxObwNvnJOPaBFo3wxSbFLSjAStIk0UVNi7JSb
hXMHCLL1IYr8NOv7QqxSubEu1M7XbVt5XhkAgdw78qWDXXCql0GqwH17+8uz4EceqFnzT4a+rxlV
NdzLDwpMJWJrC/5aF4ARCV1RrzoJJekOX8kAFjR1PkguJcaZ/HsgcInoyrbsaudipsqcU11q3bON
BpjPBa9cE0GclWTwOTK9q+Yl5HkrFowgeMq8EyST44MO89MYQKvybKNVfiIcw95MuLVa3PJ9tSTx
3/rb752QT3pHwn8OE7FGjvkcnHu1ef3fkCB9ToG3QwRU4w1OhaI1qeZMRPWOleQdGE5PFlkROlMA
qObSY4637tGBBHEjIwLTbgdZfM3i3yC1eWFwxYXKWk9Q6RcLn147Oh8sPIxiT4MSt8awwsL8eGjh
PZNN8/f4lxpK9L6Pq6QFEZARoGGqsA5Sbv9zLaw+cKbPRKACT8Z1dbb/7S4/99UeNxkl+n2V0PiP
wCoG7qDtyURdFz2YJfTlXNfQrru4v115o8yrKon9bLsu/tUGJj1ZfsCyZpQSM8yjJsQK51KpVXo1
/yztRiBP51xCh+SF55SUV+XagQtp2aNzuu02Y62uZs7mdk1S9QxvTX/0E/GC/T2PVJo51BSJ1RCE
VFUk2LQSOU8N2PFGvT8aDXFV9P6v1MoYtT/qJ53GiqOe71YDjz3ou8zIJsTcW3/WoiJtcstwCXjC
RCP1x3m5PDTaD5VtdIvSNBWuY/NSK6zhQ4ei0rwGftxUW0n1PXJOGemFwaPWAU+ugG0S1HRs1uet
vAb9jryzZ/hxU6FZP5vCQqCmt/i/CMikEA1q6X2xRT6HsJHh9Nc19poPAOAG0XFGev6AZFheJn68
5Z2HsGn9ZPL0gd6gNLLiOq6Agrb81pBZxgCjSPVMVSJysLA41Aw333FZgEKEy96zGiQ5k5ZiqYKp
SboOomPyJFIiDEjKGfkYX6N5crmu1XzMvLloyb5ktfjCzDhcnwXwdbHhVf8XYN/+Lv+d9KwEHhKM
M9LqEHpHx7VOhXDMby2Vp8Fe/YvQIqoxK98t8ujuD3rR4yg0hWFf+JOGHeheK0iEws7gtVGA8nGI
YlPZLqprKsOwpbwUwJM6fkIA55UXAGwfAl4CNzeVgBijXsVEJMDoWzpfhCkA7MORW8xd3y7oOK8e
/AOKlcXN+9TSIrmm6woWcrEt56OtLVRAmgspdXVSHObijSmwjjxPy40ZXMWMRx8NLdr75U0x8GGi
oKGH7ADeKtfGrSMEVhf1CZhoaEnv1z6tqqHfWLfgcFFIul4fHbv4Nqpo9dn8mSp10Hv+HAhf+tbd
tqW27MsX2nmzPjXvpipZKyfzrwLgvSmSxirI/z0m3jnhlgGDfDxe7h2czitj47ADod5W6l74AJUf
wzLN1Ap/7zYkvXXNXONWtJbuGYiSlEnC4oI5+JyOsqMVvS+J1ISNzW3XlQ7wq0c+OXbpxO1HURds
GbkQbNCjsKIR1H9RCLzihad1mQ3IjXo6Es7JSe2ykNnqnXToTAh6ZSS03yZ86tK1tU4wIcp1ZvMA
tUm1Tv0BnhvZm/qEbWNYkDxvoLmPp9r+klRCPmQqxN9F+UNTojw0iPVcmC5PDUO+imNgUNTwMEz8
V40nt9jJ5njoc4OSbM0ZAGHIAWVUOZLVzp3wELVEKgoMjSHWuTiQXq6vemy0JTf1D3ocZJigJyEp
FONg+qDEUuwjI6H7kc2f7gu3SLaj3TQAWMoinrICcx0UdPHkdZEr4IWCxMTF0P6FyG0YtL8EczbY
+RdpIaAmgMiESIm6iQVgqA+wovj5H2jqdwkYNVhLxOOLMrBkGS+wOfZVHw9NJB4NZC0pNiUnsntw
S7t4uNx9YK+52ENn65ETT6BxNfDGiirrrUOClNUbTGMfe3lIj5Uo1EEL1cmukw/wagXmDjg7zGZv
EUC4XKw8QeKdsBA9/Yh1pzNS+krHQRuQ7tf+D2i1SWHUPpWTc77bUYUAX6+uVf3UXl3L3OeORuHQ
eFSvZjsSg7NnWtNlDYJX1ikiPDHFPOnP8Oa6Ra0FJcGhkFvXVtdA3+ghW+exc6CrZOzsbuUMEDvn
iTdOj8UtYQVpxNHEWiuLPhng6WXjlQlzUIMEQjYaFWTQ119uNe+oL9XXh/xephdLt+LVDDdtotGH
DqFqMjZk7boqDrf8CFhTdJ3iTRsWyOYCggRuDW4Vl9e3ig9otDXRwTIZAmF6YfRR48JumjXCEJT8
Ov3rK7SejdcMeX2dJqRqOf+XhUFpdakKZslpIs0U75FjEE6DFuwLhG4cDVenIAjEufw4gsLt3pP4
PWbAAj8x6+N+Y9SpWh4ae+6LxeZBdADxvit1EEjQoPUjlFki/7sWAdjHG2wlmbVd2GzBDfRA5m78
TbHTR+OUSUn9dD7XHcWomNjI9gpXPLmN13B//usvWksP/2ezlSjxP5yHqvSaIpmUIEwJUAntlbN8
lZxZjowVsadXXU/kneFECvof4sS8Zfs3CCMe4yuc2kdcJcQ7zqLy6al0xYb83GNp3eO82UO5ILom
rh+S4ns8lotsOijtV2qa5cExViJPPVSDyAXK5anrpcNy6V0TlgjjNwz+9jODjhOSLdJc+G199MZM
y304g+iJqnHJqfc2wcpoNhAKggtiX3+PrCqKNHvhPogayHkdIkeav1sEeUXnqWjvJTPt0gCAUjHg
IsK5T2kOLcHj1NiPWzHDbY7DwKKDfVpDfd5vWtPuWqkXjD3G7u7TkER+xrHCxPOn3hucL68byMMl
JQFnxwhfA/mAftgnXuQRyNOAIIWNUbrguPHwySkdLh4KYHx931dBu/VKh8CafgTRCeEHBYHs1zoE
unLeQPvwG0ZLIhRMammoQnatB//YhYM7FAT3t0iqzVcAYysmktHFm0jdRWBL4+OCSEJyw/ihnpI1
BYXfANT3kCnW268R9QXHq/NU/a1xmqJxXuFJqNBT3zjRhzyLdhjytc5HZy/l6J3T6A/7jqNqv4T0
U2+Ze3ezEUSBtXRVWd+/+JVlwkZSXhtrZIiMaPs6YkPYr737XWWPg924x32moFjNTT/PXrNCDi39
Jpz3OUGyNmGelYvPUPm1vEZylOyivkZp/yIshocnzb5/Obgw0OnnSmkyC87avGM6dONTdn6zRU9K
lVWqXTl3ntO2U6IGWAcH1oI9s9czk9fcA6JP5Sdu4xQ0QhauTbWIqwgg4PfSPwqDD+maTMLdrCzE
w6wJummMEUtJZrOgjvDt+2YD9d1bR9dKlHgk/EyPz+Ks1fu9AOk63FKz4vh5F3C9AuU0r7C8VQiO
bNnQgubXOkDkQQCw4mxgnieNjOt/rbSVKhpJDyL6Hb7ytFahIVhGZLy12xERP6BQNpJcGzDf09w0
WxTwdh8HBP0kVKoWKmkH7ouCLsaYQVfmeCyITn7J7eUKmS9+rg4DBZ+dRu3IRmyyKEpTDirDGi+v
Gfm2a9pH+9TBRyrOh88yKA0Ie9M2drFRXc4FcUmlWLT9LF7e7VprvEYHgyqgFBeB1Vu+PvO8kkT9
cHDhw+9Q+XeJ/wuA6KW4InZ6ew/VhqvXU2cF0E2BPgyYHbmkWAjVgVaTxG6P/yqU70xTbTp/NSbN
9cMUGF8Y7KDXKtvxLvSJ/NJ7fFM0XbizS/vQoNrQ9Hv1UDhoAThOT9zMsKfc8pGNZLcaCc+mL6Az
eaSjKqeCIAQemkG5tJ1LmRoug9xX9ofr7f/aoRSJkyiDj9dgwWSEsZsCyBkEdMJtuq6PiwO/jQZ3
1bj4pHFcALdHe/r5nr6pfhBtf7VeR+JRRAFyrqrfGJkh+70AaHdj11gSqnw35j9rB1QWGwEH00E8
PX3klNqBu81+uPgb+eQHPQTxD+cI1zMmXhKBC1f2wWWrIYZMUsi+KbjzOqhraDsVwbBZ/gSxhcT8
admzK+FosGG9O02l/9NWBrnQA1gjDhU6ZZW2TJW1fAwufce+XE5oQlvA6n5mk01V1jXU87m5BYmR
FfDbmnOu0JGa786Srjqla9NNRswOnwde7fjIZ0306aAdOn04x0w1qs/Zby4rg1lB/+BbXzzjILS1
fUrkh/LLjFMlcvF/WVdyaEnomy/9FbpBhsZx/EmC0c3WnHNkmylM/f3qqX73kkow1+HxGc7I7tLr
o9sqsV47GcTER19isWpNSTj/z8UxWHJKRlow6oE+lsRyoz3ezHSEWKX8Vz4SxMI45V+MpHvIDGmP
sW4DWMh2Q5yT/yLd07o3l6SZPsSfmNZeYrWyhRcA76KGRegz3+xulEdjTrsE8TDNkxO4QnPwflXV
IuqYgUwFE4KH8ka9BFr12DISNtt1vSxYECHhC42/t4VA2bX0UoRe9rY9SkpU/kfHv6vQseygMLXS
qiiz0GmSm/LDiu0ituMjQuqTHBzS/G7wOQpSdEi9gnJTBsVafrQgnOgyC7ODxG4PnjpePQmhjKur
HgZ5t5LnElzKOdk+RHPRJiXoMnjcZ24QQXb/DJDYLevoEZurVDAHBXdhiptGIARXnjFxh3kbPlGB
h9jChrdKI7mkv/24fVKwv59hjVUr6EydTHJh8cERWiR9Bk+yKYwvWqY0wB2vBy59rkCsqqZaeN5w
InrWM/qu10DbbpziccAPENHSvJ8XtJiIye9MVMKP/kT/TzsODIVdNdD/mGAHIwhtz80AdLqKCcEq
jEqKvwz1SdpxTvGt08mHLTxKMmHdpqdkauIH4A1KAm6IpcIVaYVIFG1bAyXVnUIgelL2q4g5Yniu
XMMjMW2F50WdAQKfyBxCpmFumlTDJ7JHZCAaQy2jScmRGC/ZA32EFUeg1DA6hoH1yKfFwaZ4Jrhf
FsSiw50P71wLLr7xN4lMnEVsp0uYU5ecafng9LD1+2pdvVqrEIChAIAgQAtpS2YU8d07hpKnQJh2
PHQMGSN0jvAIlDHAvEL9xPSQlBwoCx2EtWVJESVfQQnsMgiViKzQmOvQtogXJXvJfBnQSpZfNMOy
/m6ZqoYCY3jHeLfj18l+ZYut6azd6jPmxMivdB92YgMEx3sGqxtsw9rQBRlwgyhxGUQhAvsBWUpj
2fNrc4dYXacLyUyrHgYVP3yRaqG6O/Px57FQcuoP0C8bkvdDiBcIrdmAq3Xsb8ANvMebPJ9KndRX
8zwZlftMleZg28rarm03k1E0zW+U0k6XP8gifzJBi0ul/EAEmXKU/GxNWMJ6k5RI/5ALvvMsusad
y2/P00Hp41jjHj3lo/ULuldWOdKabq8ADF3IZwLlZWr5EWkFqYAlwvJN/YAq2vY9HiXEnldPoskl
5ZmGM8w6zQuclFcVVTEuN/FjmDH093UmXgRdF3l5jRYfxaFSui1eQg9avrtDU3QqbvqjCRt7A1WX
FtJuoFP8Jp4dw7+TqD8ophME/K3XyGOmuaIbawFicszMR4iDBwVn7q5aHqlD76ReryfLS8IVLXQO
lflB6801oB+gN8T+YZxyIkOgvftcdshBs11nVZ6WDqGXDjAVy6OsoGo3LXdkEkMsa+3mjzjyQZid
gefX2wYie6wgPp1EKFvYcCq2BCqKPFZJQIFjnYFhivGrEvUBI0t3+V97+vaNNwS8u7pnU296+sFN
cVtR2+xZuJFO9Y9m8Esa21W6bq/hdCq806xv67066Y1D0wc99uAg3kq39A7t2JMyeisgOY9jXasU
gkNP9XHkG1ryaduaNd+L+XaSum2blP56dApQpSqKMJk1q0GlNj3fyLHyN0x7ZtWwkPbKbh9ZEP6g
UUyxI2DQCSipCe0RtzujQVX7Zn9YLGxckel98Eso0LjDUJVLg7Mzu12tHJkRpeG0irYHRtMBCJSj
qFSuKRxNIOXIEoXc5REKVwN1kAS8KjCnxOUEwEg09Fw/Yo827TYvf2v0o2u345gqoNPF/ktVgQS1
hcYrd6G1PswlmBaUJq1oBojX/XYi2Qiio1ThjIzNVtAYkuOd9k/17RqF1QEWd8HoBuEurgznt0nc
F+V3peX7UE+PZgJ4U/TepuAIseNs/W7LcoHMckzM2hJ9q04c4qrH0Q528gOojqNGmTuNeciTjGAe
ql/kqIMewm8K2jHromADSQAdbEbLCNODxJHkf796wtdnVRIo/plmBZsippRUCdd/7Cx0oW2eCsoW
jZzFRdyuMsC/oFMjTZspHb24pqEgyTtYrNHBMUOFXSA2vQd979NDlG5fU3aO4XEzreiGhWsNWk1t
1Y662N04a6VMDg/NH8vGiKzOsRjrhvu7XLSZPm8m+XtXwS6QhcdjTqxuJc+6wBUrJ8oORNGL0MVU
OFdzEVYTqDhP13vnINL1TpOPl1PfXBKz0DZ5/xoZTb/5AU3GOkLEmLiWFNvF1ympVvOD4v9C/Czo
Od9hffJ0GcJxosgdPsHzNosnOZ+NTx0k1oMASh4eKry+PBu4kKVe3Btdw+Hg1jFJi8Vga2miMkHt
btQ+wUVDYtWkSBJ8LknXfVsXx1t6g1pDglFeACGG3S5kyEtop/TtShoXLNuQW0xFC5XY1+hYSpst
XOq9m9C5RAfnx0wm6UqT+onY9neOO9Safsab1QilKXoMnivgTORK7mKGwzJBZggFTQhVV4Cd/lgn
+W1+/GEbuobqeKcKWNBFcwHJSgKMDseWe/pp/dd4KBcfP6Ro2Q+/1+CGEPMi4FAzT+QfOVIUTDD+
Exem+lkoTMIz+pGpAIfZkhPhI9X5tezmiJvmSwnx1+eSviqMel9WKikkEVpl+oTbyqePkAwCO81S
XjjsCZED7+skvRJG1gNGVHLBvtsaZt4rB1g5u/RVW41rP2c+cofagaOagT8OWJHdgKs0zx+if5sW
b0oZWXdHrprZabFX5npMYzR9FUmddV3G/xE0Jr/YgBCTF7SHpSSoHVxjaF6f7ntHtjJ7KaiDiE4H
9yt1oEiBRbGLAe5ciClo7tN4fTWsvKtj3CjkLzF4UpcoSUw9heL+QZelgmUW8c+CG4UPtxTkJbAi
E3tTDCA7EayaiaHQehq33oKPTfalpG00wxp05vMyIMjq7El7bTc7H01MpKlYCAHi2NPBh6l/czT9
sFC5eO0I/7ksAgkZ0B8vdMEFzafF/22ppAqSPjeMNpRsHkDpEJ7pSFx9MWeSTrSIFcM8wKQwTPdo
4Y/P4rK+3VAzFYqgmyGAz+05FKxi98uqG6OCLiQ39/sfTQga9fRGQtHN9+Xm6YLbRyInZfruzdHl
GqHZTKP0WQIekde3gb7v+WHDtNa/tLTOGlypWfJ9sFxa69DQ5OMOIKV+fSF5N0cnb23+eryoEp4y
6dXR2aZPsY2nPcIYlzdpapVlHp2iT8m3DHIG4CFuTpi/CliDjDXgv+bYOhBISgI17FLiXzOc4QXb
qAIb4INYhHLY7cZFDE88Cx1TH2681COm4pvcpV/NvXKvIktmPHx4gZmLmQ7jQyHpp2vESgAeyjLr
rpMtjmstvJuEBJDTnCK98unN4jd2+JsO3fwK50zPtVKo70O+m59C9jVKPooqbNS7jA9gyhTfCQ0B
7SZRb9t73bBUY+7aln6Q47qQZ2UqGoEdVHYz9nh2FBef0MQW/hi83tl/VJgV4qYelQfITMmzY+nX
d4wOHsiX58O5H7Q9x+R9Z+sCnZJvhLGC2dsjmBfuttQoy6BfCbV9/WXDnuY3HmpZ+e/VYbBfNIY7
cKz/m7hFRXOGR4eWGlSkuotkYdvo9rXMJU0X39k7ZDLjGdUZsSFW3yoqb81x7OtnY6WaSAcDZORA
Q0xD/SlXfZbCOc/+se2/1UjDNmCev8Z7pm4vt72Wjkiw/2I8uPHU0LQVVaZl1JWXCHtRN93qN+Hc
wJtnGvAOEY94nfDdRdrR4nTAWUSbEq07sGrEx0GI3C0LXAboUqAzuJR4jRP7Lu9Z3yFqvCnGd6MO
DD581J1G/ewYm9TSgrLMNycT892F3Eq7rjJcGIejE5/7E1PSXM+ccPA8A68X2ztyMEf/ygukLxyb
SnCru5Rtz+k6fOwzA5yV2myjT0tpJZqm5dtwC27j2PDX/J54vlrvR7JXebNTA0mVM7sP7AyeR1PM
zGkGxBosvz0iDhMlMOUTsrsP9R7AMXnE2uFsuQVDvmSCPDEbG4Ing33HmOQqysxH4XcqtatCO5CZ
FIiAwiYGA8sOEQS6GMHbY0cti6PSqymPN8pMF5sirzSmNdgfmbuOEoz/OAkMCYWBx/sp33T3mvqY
jqOzjlB54737wg+opVgfbMg0xZoQVb6z3o/TL9P18R3teBHA5yYJMvK0jbeB5xsrse47zOHjXW/X
aur0mwrQJK3Em49MVn2Lkl0eHRMx4MJfKHVpW/nP20WgUsadc44duQmMzb1lT51/+nSTgqiXLbo/
c9eMXUgQcoTSteJZZs7tUCNZ73VtYBTEsgmD483UNlpqCj/beL7AB9qrpE3FJR7QXR+2Dzaa6Q1y
yZHq20wxQ0vlneWx0cAC7Zef7dz6jv3IKjtNXI5ecZMxzFwOWFocdjPAe9Ecdp48My9hPrWV3yi3
keIhzPZqM0MZ05mqfjM84MCurWjTVrY1WoBoO3xCwQAEF4LjPOU9WnKoVYxSa5NEgLnGREn9CSmn
zLJRuy8us0+njTHnYchu6/9pcDz8Ij2CF38rsJh1QhYe/0L8zkSdST0dDY/o+SILRLE2kknfLIur
rJdznHVKeMzFbMgIMyz53ndKNK9NqPnMvFL1uaViU0KjrMg811UvFDnUeXHvjapxcPBhS8xXTw0y
A+rnSj0XIVhMnzMyJBI8fortFPGx/q/7PmRwkvIv2+eL+lt/KWyfvPMGu8M20Y6RbAaVKIeuyl9Y
GOYkOyT+3YjFWzwRPSlz76xMrUpx/lnO+yCCcwTec+y/y6rSK2UVy89VQ1g+9KRwPIDmJLK2YhAi
L0wjZCjX/GpYjVC30mkKq2MYyk4pFbAiH1ffE3D1CJenddKbdd1oqgvfSmMJBIJYYaUW9IDKlxfW
Uv25o8ae6e4LfATpPRmuYIXyRgOw69V/xCGA7AvWX0Ons6EVYFlxbNx4rfEzM+PtwffdnL5IU6OA
PNaagPVegusu964mLyhaVunWy7RTgIRlNAhteJxpuK8PzKtKOWA94YA/Um0i9w+hI4ZwwqDO9Kwn
SYZTDj+TyxWDu5Mh9b05g7ajH4ydn9WUDuiuAFcH29crr0R0bWv/BlygJ+/pFv9i6oqcKL+quWCW
e37VzyiaP9liPf0uDwS33iXIRqObTKtYoxPKWcrnMX0Rh344ItUteOxtAPw26C0NsgvBKkgKgqKp
SiPrSrHg5al9GH6wUhz0O7C/d9d3R1QkFYU5io0K4UeBS445UScRYB0RMjjzarU7WIjNnq7LcMhS
nJJxlLJSWC0DaJm4pNtyeK2qNpV0ksAqTWBDP9e+5eLe72LShqMncXRqqINiEPef2f1lJpem5hsh
H3sOqezsK0MOmEqgkEafE3Fez5GxNYSLiyYaEilhBtvPGJ367Fk30JkyrY9qJzCMPxm7CFaFfAeX
nNAU2ajneBMubLrWUz6RBvo94Uls1Hk1MeA213zXEUmYaBXNS3xbOc/FqfXMcT/3hCYZMEbMeeSt
0NZIGCXRjxm/pijy/2RjZO8I8JNRl/+qDxD6PsNwe+dXlTPM1Pc5Pw7GJv8mave2G28yCkOw1LVp
jEZq5dJhnW/xRiLS2QzhwMM6ICFW7srVqBk9ncbq0itMAWsGKTYphWn1NEuXzx+cQO67+vyr17lX
SUgx9FuOfhM0LRA3i2YoxTiGqie6MLARrUKwjT2u/Q1z/7BtQ9T0A1e7kRcFAFBd62N0hfwrrAhY
iqphDV/pJSpvcpyjRDfePqaT0Wcbjdca4FdVMiYKyKt3DepQHkQOY0yp8OOLUMBltJixVuFhxUs/
Nv0HF6EaVwvOxRoizTRD9CcTmJza0D1TZeEbmBpwegEwC5XpQuK+jk7yuni956BCeIg1RYFOLBTg
Z6EKSzz/KD58PaJuZ6pvlxBzqfVLC+zUqBy5fbwNJsSrYZ8yRJo3xIGPp9lqi5N6sLescpP1p0Bf
oHwK/xacXwnjhYgpQV54CLz+ic0rkZpnbyN6H1yMRy+dMONzOJPkk0KGQIIIdxnI9a84oCqWscSd
hp8vSULiPCekX0uemDIF4bd2lrrIAihS7cwyoqLxgUS9y3TASl8f5mC6hCGbAA36FkieFVVdBnqb
KYvfX4jEZrfJKdurGnf08thjzBlISip08mqZ0A/VuDFtrIO5u154Qcf2i/xqtaLZZHZ/Oo2oZugV
QASu8JUNxXbaVN+vYX9IGlXPTeTJSD4nv48AOTx6qsiLq+lNZyQ9yhVa++fZZ4I3YKZzvBCTeqUj
8qvUBYzfRuBaKPDA93seZQeIqqYnoTC0KYSUEbrX9s7aaxiEhZPEdYfPB//WjzW+iBCmXgv2cKYb
WjHIHusb8CQZBMdS0zvlGgPP/zdATqeXwuxbtGq+AohOTbRgf6FPVWTwOvgOwNHqskm19fHFo/pw
RVpPmXcYY30FR34T+zJdVjYlhVqkvAizcXKvACRbhg4+Ps9rpX6+tDhvNCzHpoZAr02uzWFbqNi+
I4MBHRd2eV4sKRxWGCeI0rnVAjqNMtFQ8RuG5ZgjVptUCB32oqdy7SxlOejgPtK+QcDtkpfOLzVD
XrlCAMzPGYbhcut/iKIHlhukiuevVu4+jUSDVq4JKgiUwGoEWIMN79Rtm84nTjTBKVqeB5Sn9gS7
3RV185sK/fRy2rkv/XWZlZCtfAMuveFc1Hkp6hf/8J9Zz1/yZu3kbHnO5zI70mvmus23kzJ75xuA
o0WLDwbnilDHErAo+EKSGWqQAxzEocVm29PPg42jhq5mNADi81xUHVqewqhf1ScOiAQDVZ0vfZjP
jVX9duNyooGZral4iZXy3XnOwZwy5Kgds09pVEdJkjNUucuDjvoYrAsfCZlQi002nEYka9Eq/pEr
UGHfxdB1Oe69lZn2AzjyEJZ4omOo6eIb7a4aVFPnhcT6hX4H9FOD9l1JtbCqxqMMJnQ90FGNqUqJ
tiGtdZi9Y56H/YErk2ikwdjr1Dkah+ZEV5LLIyp3Qt3tqRTRHFjBILYY+mjKXc3Bw67aiwq1py+5
UbKhMCWkYV8wXyn861QHr3Ulh1EBERZD7Pwwb/CMXMWIAwFCaIU2KtQyxzlbySwUoR9hCvmiFWmm
Ssnuy628HpFnGcX55I99hELNncV6yfW2Wd5xQAZQyz+r8b+oDHq7O3V7Wz0Fl+iHJRvL65Nck78q
WPL9qoP+pjL9wPWxMEzTN2StFgNxx/ucDjQEq1Y6QnG2DTNWppvFf65YqnBMhlNwdIDJrTJEukeS
HmKItfiRXvV5uXVBZTS5KqkJx0nhswTNSwm/Q11R9TWbn+9JmlVg4nDAOxBJTzSO9xxQBVVcSJPv
pUnnOUN8ZMwJmLM27QKC7tHSWptcjuBYbuJufWSghBLpOXpnDAraYcIHvzSzdBeAIa1YDBqPE7np
rIrLA0qXHXydbH6wb2ua23Rf6t/DPLVK94+L1PmDuEqyyi2uZGFxdJnXxLTae38gyfMTq93GVoTN
5AXw4h8UnCeZU0F78uz4ygDbXayl0SH7lAoB1vhvZDARJhylbX7H5cClJO4tq8nA9cH3Up8rf2+w
MzgGhiTGDmM4obK0MRjgpJQvz1IdnQdSTh14uqqeuTvZEZR7bMOrwZtwf6Uvy4gLvXMS1g159Hki
zDfQkMmj0J0AFS+7nXjX72iDL3Nqc1usSuQ+Gc6ItGRyh+Kd9dXvgboZxbgiTzeBrfnQZRRBH9rh
MQkvJs0fuXt7/PgxKFN/qR6WgGrr21O9nfR0JxY9dXK+IGbvcocVr+KS5G/voLUxgHWOG5Y2T5q7
SLOBMXUYxmQiniYsmAOy90qLkZRMbCI+1FYuFUKpSiwd2aL8aiQuNGypUi8l0JGd7uVQcfnGmwzB
8GVmo7+hTCIUigy4gAyn0c+ZF8FZkk3EhbJFbpGJBi+gZYpLScM2nxed+eKingrm5j6BLsP0QS3b
GwuQXpGDtn18wULIoK7yiG/MNCm4Cs9VR9vtbd0iM19OYT/FhsDVQgm3GIvFy5nkfojejCM71lxu
fsiXESnobkwfKiUoIWd4p9itbvxGWaRTXsOPRPVW5NfFmh9BSbr2gUHGNS0lCz7q0E3lF+0g6fXj
gEEbly8XuFMGm9mEwFR6NIsWbe3HLUxprFaJGfdMsof9IhX4cMJtg/qv+2k6upuAOX3p5gofjrH5
bHrwtgP25KgrZZHO3hMKAtTuRPmoe2NyC7+xRMGJF+bm7wQFBXX1yUvuzI9raMdGe3AC7dCiw/qB
6ezQZcx4UqL5tsbVFvkyrd1vX7IF7FNRaZEBguRtPdkFggzlS6IJcvG8o3tWliO7yrJ3AREPeCSC
Q642Nj4gycVXUpy3K9NtpZ+e1jetxULMC/Lzsy6c1lpx1lXxhfyZ2MVdgz1fYuXJe527Wt9O0OKn
2Ky2r7tcYyRneCE/jl0gnq5xf5+xPPigBC1sp7tDnI2+xEx4MaCwWZkkkdKHuFJip19OKC5NFF+Y
PWKSaxFCPQm274Ok+TjK5djrj8cQd6Ea95WuXiUiNPmNgYiFSqMvVjTAjwvhfidCHzZKBUlEQPo/
Mun/zQhFVLNOl/rKo6rt3ixu4HUBsBWhs/x2h+ceY4LI4BgpdNXqr543OPbb5Te6Mhuv4YtKOR9U
+XUkbvSPzhs0ulL2uqw5tRNySUYAxeytIwpSTgEH9N4lHgBIC8gbZGIY+dXY4wCm6UU88aBi06mT
9NZHTuwa6v5QbiFIfIYbREVn5TbM02qI88V7QMBUHHyY2QuWBPLHJ0PG+lDmA98ab0caPbAIXLCU
apKmhEuXAVXQ+xeKcLPJypArEcKiJwBNbANNnPXwTUsnj/V33W3t9GX914wtyZYUxkenmNnEltrA
/sZpBQNtsStw2620dLi/xQ8+YCSuepIPY1WqGJeNQnBUvsMuDzNjkTGfpRlONRwtr46KETb3D84M
BkmoGX6p5hFQ4Mtqxt7ZVgOVJ7+AOOKABfBP/A/K+K5APF57kHkLPK85KJzC+ylfTNYt0F3oe/cn
PChIJiw4W8B3wICmTNPIMZylqp0iGmFuGlCzRweSRR/Q9vNpOCKQqAyQDy8Tf9aCqSFkO2xNTV7m
6anLSk1550ZAO51oZdWofqdcqfCbMg8SZV5q2GXW+Ag/FVv+erZIiWIZ9+R9HeQlAwZ3zGA7qdrL
GseZFX7hkdhSouxjbh+YPPOHbIWLl6vAaEGV1a89OwP8NkHrt63gNsracX8pQ+uJ6wAGtz5gNs8L
szId0IgPqUbJho5Gx4kIm0IMSni9/EpxqBCkV3JGohcaV0KR+GX+kKAQ3MF4MaaVaTq6XidId3So
GKTAUFHL5Tksn8dyHSeKzwFdUkkvdBLgMzVQNscTk79QLFjUUtdzO+cSJR47RuJe8+vlOBVPRRUu
cfNl8ZjXgDz56vVHT0aWJZ0c14JlpmF9Zl7l5zRJLBlPg38lIpQpQAoLvsmG2c/scl1tMMNWCjfC
9jaJoHIvXGWVU0B5JSdtiZtGalQLsrRlmWH+GAiJ1DlILxSdemVgIqEfsWKIQr2BN2feH4rXW8SL
j2heS2BF+BcoWZDiDfxHqxZYq7DsOfWIPQTvcysj8P3D6FVyeghHwyIYMw4tJMnvBoU5RhvoDNS1
r3q1kJ6i6XjXemaamgVfgfOS5W+ulvajLrr4jn8T35xLzo+IBQtQTJc8mPjyLoCWMXI33iofRbt/
E4dKzTFHZaRb801gW2qsS2g+KEunTtxRyXVDW8NQE6Vp/UyjJ96U/Ggs39wm7Bib1jVjNiMMYHx3
v55e8GyQdEE2N+eHMGm+NLDUAyDLy9Y9VopTnZyG98KwhRddQchW/EE1Los53xNP4mv0thQJ83Ca
kSE8gBOGYtkGaWayhLVtk4W14ublPRmdg+PVUJvBw/FMT41WsZ3hJHcuHkLYX8YimtECWz4whtBe
g4bMoXZK2SjqYJzcKSaDUckfMNhOGPF/UUooOeKLC/Hg67WqCWDSdzpNyL+KBeW3eIVKrKQjtld0
ZYmLHjcDuXX6ssBNIWocBjw5fwrWo55LhnM4YcCHpx7BVuhI2+7tV30Bc4Lm2YNOt5uW6ZrMnKLY
+MNZiPDVjp7gG9pfg88qSx+GKKFTWYUTiD/v5kKsP0HSNroVFM0nBEJW6G7KPp/QrbEbGb/Ld60X
JIRI2ZGl8LySJ197q9SzMqmiyWkA7n/2MDGAV+yO/rfr7gPEhFUhYQv/dYGtBNyS7f2m8Z4K0Nva
8Noed0+wydgkdBhl6ZsMlm6onsjO7v2DeWmiSrn5toBpwxrstp1w8YKXcP2a6EiDPj9n07B/NFKs
0iJYNPCqMjclS8Co54acg5rSfbO7ZfZRX1F6Tlm5fmH1zKlEn2oSIBW2bK5H9vILq/I1+5h4D6ie
OoS1RODf8sfoKSuavWz2Gkod8p9HugUYzegJxjTKj7hWfU1mK9Jtoy+OFkol5A5wmofW2Y/dUzhH
nB5RJtD7mvPlh8CZgMzqzPM0Pl+Y6yLOoW5gt4rJhso8LW7exrHQHe7UPOB8D9Q4LVpk9Y7/M+o2
U8lLzch5ThL/WtGnFxz4CIx6QbB5GhVYyIh8dnfiH8x5WpoiRw/KkA89rGSaRDl4aqH8ACgwr3nj
qC/bPrnVMtS0bvnuvIVbBc8cbcFmZ96ozcZzdscvyn5eAEzNaSrhbCdDgn1wYvf/wOu+P+51HRmo
ir54TCJiNdxZ+Rn9/ycSuP8VjJXOIgYpgSMHMEQ+EKUcpwwv/9GXr5X6s+D9wVe/J7hbzRyqpOS1
bKvvZR3TgqXS46Rdk6n25J0XkZi1MschJ1mNFVvgVutS3W1OmjiCjEFGTOkOj21/0nPAjod5Djvj
7+z255nbxj6S+8OqgudQ+OyC83EAsOYBorJk0FljbDOqmbFRwr62P0AvcRKgyxAU67CDEZXnrlLd
6kjQj0uhETlFbRWKrmY9Zq16vLOFkHdv7LojreAKJIXuBcE+YTbSDXkpJH77x/CfPvFxxlUhxklj
YxdUSyVd13ksKTQ7D3yumhswD08n05FBBkOyk4NCmy48BeW74FkPK1n49igrCeMfo6mzzHOXs2vi
wsJkKPq5r158LC4Tyx20CnFSGBAZ0/LKIQn+VDNwjX+L+25gI1bJPUK35u5oWNP2T8636CA9sgCT
mq7O1w2VSAFdfSqpZhY2zaIbu2oVTBNiy0boHUkpewOs7FvAlSPnk+u3+XWdAQ+BNCuVbHqKR+BL
kiE7pAQos9SeBhWzvdFCVmvU5IjRUmdZRozzFG+gKd4oSRg0P0G3YUyfkQ9XZHmQqe28ch3shp5J
YnTstXc2uXGgc1r6mYugxVyVOjPKBOo9OCMJyxqxfiihgLxHeEpnaIKeG9z8g+BPf0GioloxdjRm
GoZI5TDgrZgEbpH0v5PaMj5xxDsDDZb0CukBC4BFql3IuoJldMHfjC/MNZVBCHa1eGig8AwXna+9
u4a+QvffpnJEzH8fRYh6lM9VEXk8AaYy0gWrTEurPBpkwBwqJpw/jzLRACaeeCasxoZyoUyl2qXN
n3x+mlA5aYF9CDvMzOcjoePZQL82byV7tXVQZNC7FqGmcKGEMBo/1Ymj2DLZfs0vzspsqjqrMrJe
c+P8FkhzGzJAF4ai4zJWj5LPmnGStss/puhooReWrET8N6wAl+Xz79C04IceqSWaI98NfNkw5buv
QBYTSX8yb5pTufuX+n5QG9W7NQxWOGZ7VKsqRVQsNcYo2/NApodVVwTaaf6I6PIivl65VLjKZTgS
ail01Sksqjb2FOEux+jbzM6gMuYNRiI1kcelADeVn0o2oYUPKsB2QjmLszT0N/nf2IpKjEnQabhH
V0h8lAYFM4b27BL7chY855ztLhRwFPUOR9Vaknau/flzTFrmaIkf9ou8O8Ta5vhduEJ55wLYHj0g
UqJzqp1WBY+jGKcjpzdr7kspNa+WL8aJU6GZaRyWu1xhn+sM1nSLkPr1SXckLLXyWr3wTuaaHVy7
2o7axMms74GNlm7st9BNiQf8+7T3u7xWIV/EL5UyUEebPSbuAe6uCtTtmqsrg/g5Pp50LtM74mYx
lpYJyIHGzBH7Qjdv8K/iKw+aV0RXyFVUiNnvo1SUqffk8rB6d65yDtu/z/tXg7i3mRVgFuuZGdwA
mOxFhX9k6xFYYVOJAzB3ooOVrpSO81dO6xit0vGy9cFU9DCw6w2hJIs4tpwSuujLJVfTkaPe3nVY
vWp6nFkbHDJODzG9rI1COgf6LH1D1PKe7Dr0DnjMYywJ4TQU/PUccYE5ohgY4Ka5TtgaFcTun3ZM
HYMlpqP5G07EMlOLsjMHxQGzzF2LGVpyAPTb7tTConwL8iGFZQzSmEmVnWqFi6X06wSisjpqROoN
hlC2cGpsagXuThCiu/Gy8qfk0hWF5nbaHJF7W0Pih6vKZowSt6F2gvDK9mp6nPHUBLQbVu8BSQSO
sc9SWg3mnOFHJwGrhUrE4zbb4gL6oLtxFXuUo580KaB/Y4K5LTt/LSbocBPDsTRg4v9klv44tnlR
4QpVimKOUEOkNLSM/nkRA1V3wn4VABRutfX65RvfrnZCJU5JrdYNKsmSTMWsFxpfcchjV/l2ilqR
FiCc/Lb5ruP1NLf9WDPh+Ahm4fju9RCQfqYtWuNc76DpflzggXeVD6wCoXrxrAZ9XNTeQuTIhvPd
ziD7C3R5jSkNC2+JTD6VpaPPOoRNXP4aJSIKoe2Qupvdj98rxSBSxXxzROHBZ1TnqHGxDrO2Zbua
3dCqZaWiSaeaIMCuEjoqTVN0gqEDQtWQyO4VMDf8BOjLzBq0c4KLWY63XmisGtnSkN6C8CVrEjtA
NWq6j0GzCEC7M/zInEkFoh66ZP2J5FmZdxUqDYcaDRbiheeV/e0vzW1RUSRVBWhVY9MybYsgEvDk
gxHL5HV/xmAftnhshQknbmliskC93+l7GGcBGMRs7fzGyRe8Ix5tIJfvhZYSfgK9BsdeUFlA/vFO
WFxNl2/nfkKfRolHtGoMSl9BUXh7RJg4Jn5Bc0gh7HKWKlWz5IPo1vAH+FGg4BZDc5TBdFRC9uJU
aFYbtZO9NROOH7eHH+1QPJDMTRvtD6pr+6HrLnJ+Is0QRZcUqHfI+2LlarYzjORR/erEUziV3DMm
51pj+Fmf4OGLHUVse+PUQfsRN78u9um5UiYuts2d8YPEx98nLzZcIZTeVVyT3ip7kXgugghA9cfy
6iLQplNRgxSEgq0jS6bwN8U3fO9EFw+ieapwaQTy2crNzoMfz67oDsGVwQlNB9z/OZCEhFVPoGS6
CaSgX+PLdxzNR405G9qPx/JEZYFJRHyKL+T02u4KBNYMWWrqGGu9VY2ir09PWm7eFID2SjSIKrIP
cxNUcayqoNfTr+qWcLo0QNEKGA7hd45TPCEmZQ4iCjn9PWTkwccCOWg5gYgzEjNhu6wwIRVA/yPN
bXx6rV+dTkEOxAZd0IIR4V4uXKof/+61eALHzoLPZcKEso/D3uZhOQYt++uoi2azAkyHJHFEnEd6
cANmuIPGsJoDfhhlo5/4hTvmaNY3/62CBaAJ2Y6JsaWGOV+LYd68JHUSrlPxYCJjLytew2KoV4oH
+9HwOMKAipXbBmeMu6rpFfxHa8s3zi4ss4T4cp90U+MwxB7Efn9AvaYfVgLavx8OkPK6pi4M5zer
yy/dqgRWUue5dJnATigIIa6bFij2TVz8SAxdXWEBxB+yXjfKl8sW0/ITklMOryt9xUGDOCV5725Y
BiUhldhw/rHfsZa6+Woz5fom9RFIP4E8ZuAtqPPeR215kOe6IpRQNzzkqjOf9i2ddtUwG6D3DnvD
p3esAsjzaQxuR2iQrTgMvGYVQKLHieslepxb+uL6SNNUNOMBg4rs4plltS02bvhHzFv0/c2crTex
eyht91tO43/RavdqTnjKrjSmHFJXuEc5YoW4XwdA+iZo9+yjcMHphqEJ+vzMT84bZEu5P3NZq2X7
2DRgcW3KXFGiQJTyycvblnf/u6x9Ji58YCMpYY87SL3+nzzULqsnWdUqJhFno9mx4G4EOcDDMEfN
MGIN5PgbhcWhRChjwNljIutpFn7LnwCvJscAKIUdLhMxnlfhuTCkqyd4/HWYsII3NSUuqnOZOIhI
dTRTAvgqGmXQDKGZJr7vrwUE8mdoncBFAr7dwQ8zMT+An4KNCcRQ5z5+Apn7uH18uQiQgYDtCjny
KPBrclW4wSUdu0IcRJGAYX+zvU5Nr1jpbjiZBC6ZH5N/v2wo1vNr9p09xe4xMVuO7nMFfns648/K
rC9SyK9zPB+i4SDyqQsyqmNkGFFAqeuW3N/IGHYNpA/Sbt23IF8bhWPTfvCdOHvJQNaPtj7JiUi/
21FlIsjde8fOsT5ZKL4uGPrKF7VH45+gI/iA/TMTgluoT19K1NwkX2213I1Rwfnh64ssnk3myqSX
F8JS4uHpZWWqsRxtkpHcoNvyA5KW7g8Dva7s227naRgyPXvCjeXKbzqKRO6KHTJwaAkPy6+j+0ff
Olw5tADHzZOZyKn6bTfPFdbY6Hk0K1N7Cih0E0lpxH9Av64cf9UuM/f/+axE2L04q2RKRnIXgEV4
mVDMcmR9mF7ZZMvMAFcywhIuLebXeNWSrYGapRDnUnqxzsNk5+M1rR6MPhtJR2gML44iqBy7lj40
Dq8NoYTw/mE3MOED5vbn3nViMz0zFX9Ho/XcaPlNvQ1NQ+gatkxWFGxmOm9XDNPADMGAOPjdvHgS
TVOsTg79+fStC5GwtSdFoJ8KaAu4kWEXuek5tmq2uHoIHK5uD63aQuEnX3k08moHlOPiLoNAuLtm
WHkNAYuR1aHrnxPlGzsPlfiVMl0p+yII8VuwcewnN/F+tTA1z5W+wGiaVKqg9a+1f6Imz0Ayi6Ax
9y4amx3pOLhMbdaaBFsbNv0yc5+kdOCRO+Iz79Fj+ozSB/AMUYt7ne/J0UBKuz9wx7gkbUb9G/GD
Rd40NtMzAsbL//PYOARsGTtsruSLPMfhQvKjlbm/ECkdZj7MuIxRKVrBI+jGCeZXg8v8c9ubiEQD
/G2eGuoTelooc7qiMWxE4HlcTd5u4KHfvq2DeX9C3hkZYekpllmhtRk4PVkgSL/DkSjlgbDpdB4g
9qTRfqh35Wl0KvBLTxECAbsTx7nj/xqzI9Ofy1HD6cluablKtgGrZ9JBk+ZrM+cpp/yG61xg2Ucw
Ix0FJHg9mUq/eLDl3sFPGf91BEYZQdy3FLQzR8W7ARGvVSITAWEBqPzkY5tfczQFwXbcgZUzU0kQ
NYDP4elxmET9Y4Ha5rUEQAQs9wZbiZUMtD+bAP3ShQV+6gn2CtHVt1c0iTMZAspfEhlDuKCK7+Ye
5TLU4mA26bZjwnFrkB3kml3xLCXydHDI0DhprtUV9zdwRLWcqjU047ksUDiZ+mZKTJXmPSM2mLsV
7Rb+6mLOP1ggQ9kX5MvwTiqzRmIiCIFdM9diIJvIq2tsrTtklUR0pc8TaiSoyjUPXyEBmACFKj3/
nNgthNyQpIwuzJjpf3YaACZ7c57qB+x2ax+aKqk4OJfDISLSfNYfYHTtGoN+D5Me25R8x9pGEMjI
ePCvp44KaKd420/hIM+FTDVfuiDpErHOGHsCkR0HocdOd1haJsvYxTijt/MielVk/aPoJgMiQ/yS
+Il54NMbXmIa1oWVQwzuOP3IdQCAusCHPIRKtA86leM5k82yjMtgrY/XFnG3SAV3RNjUrpJTFWmC
lVeVpGdh0jRTmoY+qB+x2hkaHT8VdTTf/B9sBoJJqQnEnReiCMyLR45zENIpKvxfMOjXEwigL4r9
eNzAxYwwKLlC/ECMwOZFxH3WEqWP3HHKvXNfxV0ftOHiDEV2YybRktdcpJRaySlD8U+6wGpziwwi
tcTlpEBAdfWo7W0+GLqgDdoJhkLPDpnN2kRFWQ8QyPnUM1vBk8vhZWmYGWsPur4eGGqIE2O+HJHu
L4954YMr42h4m41FWjAtHsLtACvokhsJujmE6watt/LUzCza6Qe1EvhQcEnKqd3QQNCOf2shLU8z
RjsE1rrBoxdaLlBkzqmCZK7H5Kaq6eq1EP93oUMueK6ijdzigDHtFra7ktda9Ws2xLY4/1loAkO+
T+bx6vJDy4lUo3PJi2gJT8fv8Fs/JndKYPCIdCwsQiIRqvAIZb1CCThYGzcFfONdyX+Vu80F7xuH
VtHHC/WQ3xxFz3gt3k/1FNH75HZN7yGRHSgTgIBw/rDnb+g4AxjhHcxq0B4lZmhDQCgH6iG50Owg
sbGRYD8ECfVK2Z521ob1/TvbyCxQ5jQscpj/BjtRtrnoIqsb82E7TCL2a1twKBFUju4uVP3PTJqp
siAq9lAYlOHEjFc9TmJ3zU71hOJU5PmPBHwNR8DbEB1MyQhohgaCRqfs2kj44dBvMPjpClE+hnrL
a8tiGLASQIg3ZGxdm4JXhV/aoJinaszI5Amby2cgDQjxs4doO9IuTPLMhvqwbk06BRtS5TjK0ULP
dMswjIZIALlIKRcLc7sYhWQ/CsVWNVZo6twnT/5eLyi84M8wkLcf6vKzrjkYGEtuslxDfHJuMtNH
t+KhWBq/IeJRDR+NEyZoavb29HC+JqRyUK3eQXFfssb2bUFFx97mHvSIEnmlE+Yf1q8IqVvrHYQz
x45Lgit/3wBW1SHnErHhKjGfIp3nrzUyQd+eygG2OBR4oBtaStxvARz8Pi0G1Wv2sSDPR/GxpXV4
yIocC0gI7kKos9sM9VVIle7M/oo3fkKqoAqu5Edb0pKem9clzj4cg0Yl4+bAXySPk+H1WZLrjBrF
iVtHbyVe/JY8M0y0KVKvCOQpvJljoCnroEoswzhvtylkEAvE7SK/98Rc+rzLYJ2/aNiosmsK7Gul
TAM/7l/9SDYBCBx17HS5Qnr2dcxC34uEq/vC0hLe+Mdq9YAIy2IesZd2OYq1RjcHdrwU6uuyPcJj
v0eSnalPYSvHB3iEzlWKLNx/VI7nGcpBAKx4ypMPFnvzz6NArNjRAuYGSCQtL1zVxKH848e65zmf
0Ad/ybvlhX078kO0ZDFuB0NGxhwbQW4OrXab/wucJqGmd2rqTTblYq9fQp6/r2ZL4nzLvaswAlIY
gsq4hNhfrvdAT9V8JEFx80YHi5JzERV+pY+CPVzAXidLitBakZTLO4B7YcHj97hJwcVR4EnHny8V
2ztCskwFNb/Ah+Smr1vS3bSPH9Y/vG8gbg9ot/snRT8+Ih7Jl60GMalGQcc+7Lz1LUdt7AJaITzX
3fwqrWsUZMpHYV2qZr/XQnneC/+upmkX3mzQ5P/UUkLrWyMJ0io3R5E1HfNQB9KU26yLyl0w5DiV
4yZv0f5czEa600FqHwDHlqsqYc6530MwSGqkupwzqgLrgh9PnlPc8p6pLFz3Sw/z4XOu8H2BHoAO
//+Y/xS+O+/YDGGaAjIlpOZa0Tn2Ii4N8xsLjx3agkPm33eV4G9NEZAODduCaVjqoEM0LH3ZNH6r
ZR5z1f2uImtnjRHOAUZR/XAPlRs8zem2dhtZ2Se66H/UwV+dhT4mbqeqDBwwlvw/x3bAHDffilRm
TkqM102MnsFJuuRgp9TNJp2ZPVx6p9+SnonuIgVYlwDwaRLgPe+7VkvUf83mjQanyvsEd77mIZMd
SLAHWq9a3WYh2/HMnfmbhr12tyBJqFPyug/Pr1D/C0/P/YXlRb2q3c7XI3lJ20VAGRkxDsw5IWp4
GX77NRzrL/DmFOb/YrIEmbZ2A1xEV5Jd6XlcSu+xfcsQvoS18lmMDRs4GdOEJ6BAT6y1Nr64ycLP
JQscGfqG9ZspeUIXbi1s2f/00EAo4LWNcpelXmdW+6kj8DLB8BCaPDlkbQjt82NlzLAwWeCCv5kH
g+HyHH1A5zYYmYfGoJkP86zmG9aAqylM2M48M8rAwNpW0lWBKg4tyHtXY1i40fuLn4w7GZpqAYuz
TGyPyU004IvbRz1aoD0s3COYE2nLr+byoBqmRfPFE4lmggS9H80JFjkJEqqJVf2uKTIrONhBtN1G
JZdn2Jp3U+qsfAc4rr6EWXBfkjmKOTkYMnSITHziIeVXW+c2JSOQT+55KMwCOQt+3cvW9Js+RDWy
EmDjxp64HBODSGJW0TvQqhpJXrqpRix8Sa5UBDBdsABGsRnIyS8byBB6nvBPujmCHOfwx5lU+0YQ
7hBSoqXJgXCWQfRXp0+VCwxsvRZM4g+tHipmNlFwlRrbJ+C0E93KNcpRm300jXGMVYT/c7ZeND4A
YX88YKYn4jNGYiRgyDi7wfPZq/mqwBbULLKn51Hm+YgmeNGoRThEpEjBGnnLQjihPFNHu2m6g2vK
R3k+EA5zePMNhNSPvuX+5t+fTf0dS4ueterXwSGWPpAazywXexNAQaf6jmqZPlnjCo4hSrk4bHTq
8kNTxGDGoFWMSPW8qp8Gm0jhgZOVwqZAkhAext0sd1y9mNEGs7R+pceEegYQ2Q3NDVrwht0X7oPb
3NV2MbQWowpOyP89+zKkY5Gvba1GaMfjBFr/7GU/02UkbJhO1KcwXDfwvnDUbz7UJJHT0lBX/I7a
+ZudeuBhorNG7Wvf3RVAoo4qmZtK00jPBLnQ76jNJcD6UqZRDDqZjKILNhnyU9+O0T2mwUGNSy8E
KrNLJKGx/mzHWVEhKjlaWeGMCXE36C+Xyb+gUZqiNMuaXAq015e40lPaaagHTrPTnueAaJ2SBqst
jd05zsrKcm0eyR0r8oTjBuJnxPP/dbDS4bzcfl3D4OdGY4MuW2Ek7Wb8OLScmf23ui/7rya9/XYq
YK3Zs5xAdqZcD8GjSaYhyAvqFxiSPLf1YLMptR829RPP+LkINYK5Fm7ZCtWzpDE3h/U35K+iMats
OoGl510hoxXCdu/lymnHgpGYiQc5ZsX5SDNMK8denbwQTzck5OpM8ejyhZWw5/b6Th5c4sRmjTrF
Nv2a7vJ9pyqw6X0XRZV40P6PGrDmg8hPT9gkSzqPZksMkU9a6kZlUwJNRfodlPDR3myTJxtM/Zfj
hfgtBL+jFANgxeMB0n0gwUiyBVqWW/Sw5zcM6G1AHVJ4j9vJGsUW4K+cab2SQ/1i77neoorvisnz
XNDLSLi707cdsERb3js6+8zSyDZgzQwRZZLOm+8T8RnA8UMot2xsRiybgz47x81WzzoyD9UC9F34
MEzcoqu6vEh/IfCC527WvDagmtpHFHGcRHEdC6sriYaYB/PNJh/CjtPBXu3vYTWGEL7+kMBRJBt7
53zHUSPhI8wycUv8Yfoq1cQDUDFciVHDlTNJCy/sptnpOyXIcfXDgpCGz/isqQzrsiOr0XLZaoOq
IwjmiYq9MR4BRb4DcBVbFk33oqeQziDMYBqrZsoHjT2ZiiRlclRHz+kaTZs9Cjp2j9hoH9vibjbJ
CsrD9YeC54st4qEeTlj11fqAo2AN4OvBRWF+z5JYc88Q61GJ9beO+3FbSTHF9uYNLrGp78Hnj+xY
jqz3MnUEFx/LjsDXaiQEc9on24f+FMqgRVn2SlNRIwWQDSBjewqtcYNDt1yTA5AvSp86RM+CueEw
sf9kkCTv2XA85h6sH9sxZWf2tNCLRV/cYt6EZOHgvQSXmxaEJvo29zBOeYWdK1eWgk/auI9tK8D8
Jq3NVy/jW8Vecme7djh0X2i+kZZy3Z4R/WqHKZdVI6Exg9s39/PTd4Nca+SJKFNQr7kvWbojdgju
fuZRPpMNRdqOSuR9w8D7hnin4d7vu+PEtHakaLoAPS8ix7XqRqrwUCSG5lsH2FRnFHI7PrghEQx7
mYEsNixV8amg+BmvVpLZZ2M1vI8uJU3v4YIbQCKeeSbo8QljxSGCyzEf7FxyjbaOsfjAetn2sZvx
1ztwZC4LhxhsJjo12bl9VEk9Q/591FSrDvjY4S9SxUTIkQtq1jVKvQv1/ivyYVSdSM2+GUztqqaM
WE51YqPQmIa4HFkbLgObkvmhwWja29Yf9aoqQ6Xa5QlwT3LRHl3eL40zZDC0GgR7JhcDVPwrOCJw
DZQNzaD1lHtINHwn35XxRSURUia74qYkEKf2W2vVZGstEyeYie8rWJUyiOBxSVsOo6/LWoeqTdqt
4mvL5L+KoGHcClS+H438sK/UCQXWUES1mQvzwyGX4VncjX+qPPr8Dgsfa6Svy7+WQ2QYBskyLJea
kRQDlLvvQTA2C6oUYfQdVoqam/07x1yaCt7BOHl/czxp9qtH64T29IJjzsuOeZ86mJ0S7Yca3t03
lsYtbQvtcYEjhhoHftlx8kC/3jbmSCT8kB2s9/xeEWr59KhnyzMvTPeMwujb9UccHG6Y46vEaFdE
DFkCHAFPN2h12r9q6vk2OqBLhWTK7WkFxj8X+R8t+2gVPGkFZTUc5i7KP2eq6xzLzC1FuAWxxx+K
fVwwTFUB7V/BuXCHwro5d77/NuGDXoRLVIm0u7IpJiWnOg60JfNbY9u6eIcL3LvnyEnwIbSDKJTT
QsSno3seUB/6JJzj+CTN07wqaqSjdjtyF2zSg3QFSgG9naHgi4dKzN2PT6Iercrp2d10w81fpDyu
udoI1S8fI+oI3df8LwddTrT/bdqG8/HsRs5sYdFC+xrIpIkzejCJNRImQqIQhOAYqONyOjRLJge0
01ce8KLByROysM3VuqAcrJ8GgZbtLBoYIl5/XeXfaMQ51rM6lfC5A0RVy/KiWTJXtr2MNUCdNHF7
5Iz80XrhMSUPAisBcjIURe6lrXKFpY3Sl4lUral9buCAylwPJt2BgjQhlFeZlaK6D8a7hCF9HKZ8
NlqG8uEIPlgLnjn6qoTtXAx7ZG9TeD79Rf7blODovfIv6E0HdC1pH1AKY2iIQcrUIBnKGdNOd1PB
xvg8y+6I9U1Ms2LrouYyIj3vQXkcgsXhXU0nnhZ1v1UXVO0JfRl7gJzjTw8HcTxbK6tL743dbWmp
gpH7/SXAJnXJZ/UHm5B/1HWe+0Q/eJr41PmC7CkjACgopeQKOprkZRQLjT6GCDYlEcx6KCYDPx5r
jtOElBcCxAYrVMHNdWqBh0NoY/8z0jpwcGZr6HAl9zwnsUiKqy19d0v9J6N/kDceTbT7wGwOtSFq
HHboFzl8c2AV5yuUbOd/HllDKO73Le8ORnjxfvmqTjLwFGh8dBrPrNSqP1S1S65jOeQZzcxmV9ex
JIwL8ZCbAEQhq/KBZz4B0tDUxKOwpUp118GLzMb59ujvyvIrYcPlMvkhkPi4+ji4C9rrHolMmEF0
4BaIcOzmkirSwouWDDf5aUF1W55zadmrKsOZ2twyRSeVN11yzOEmdyZaq/khLI4aZ6VcgNaPWMYU
TxA36xUY0WbYqunNryRk5Ez52YkgZSgg7GCYMQQeZ9Q3Qz2W3vyVYrMZ89g7l+vbEIbJ14Z3Vp8K
x0PHw4SKtxufn2s4V0GMCcYcAd9M5lhedcs3ziG8DBeSJQItwMf6NXiKyGx91sPm8/lN9dlr9kSR
LVM9yqc3Jv784g6VH888UqghhaDgT2XarfW+kvyYSUh91hhapk04FeC0qLVpqN9fqTL1s8nH4S8Z
EMV8SEBjRLtBWQumCuWalmijqErCVFTNEiG5R2PuGFsGS5kQIsPhhD3i90yfWh4cERxt2Dcaf1sH
8wTknpR9EPBnA1ncQNsNttR/fSKjRkdsVrwj+M8to3QtJwtyT9TwveYD7I38LRSwiAPbixP4mGBG
WdWrSavOY59iRb3oTQz5LmS2OgZTnjM+zqs/N6TD3c6oVD9dhtuX1AAn2EN33qx/zUf7mhe9YCcP
4H/tkS8zk5E2v8tTjh79Aiu5PjeimlJbPIMXHjyHYExQ6fjHH+x794uh+s5rf8T/PMTQtPTxBsYW
Llmv9N5cdNZF1N/F9fHms6dGa0E6brn+qCRErUStSjCCq6alIzVa4WWatg8cso1a7Mmqe3Ks/kk6
X2U81Lnu4vd4OCiStp2AMZ677EP4dlFRSMBND2SetpWJefHuRluO13d5SjCqJ/cMnp+bOH3ol/kd
ldMO0cnp/yDsV5YmUmRU2Sz95sZZNCwYvHTkR2QMfQC4ryyX5G2vGlBfIx3hw1MZ100RgL7p7yNu
c4ZOdhPHGLkb6f+O3Ojt6HMfhSHMXKdOLqDdlQT9Tm8VlkN4q4JTsyX33wY1ilUOb2bnFtmaoM5o
gm5wPVGP8kFh6aQrvUKKcCArySnTNB/RRNU2uP94woD5LEgJfh52DfLcEGowSzpcDHxPHCNFnDrI
NsbSwP/PcQqLogvDxEQdZmpHLjewIzxoCzPUX3Tli0p4CxLJ5q42h/vyS08F/BuO7jMlDesRomg1
JCCf54Ki2WlSRv9KfHjEdkBJPnGOjwvwTuxGm82yUSBoZAfnYYbDmaRT5cUJYpBpTx0UcBzK0hF3
vJ44DjkLAm9l4ciaSY3qiR+YJHg8lTC71RQIVUEWrdmLnIjptqeNEkUGABf6xzblEZK9+UYMtOou
aJ0GlX/n1FrR/J/gyHm1Xy1Svp32YR19G9uL0Fb5kr8wdcbdRjsKfBqDvcQqv90QXfy17q2kw4UN
wl2waUVVuJzQ0U8o5LcDZsOxwyUhQioTQbzx7///hjQD6SPr19AuybmkexRiJLyYR79AxKIxUewM
9zsB36fWSd1W6cvQ3Vr82WYo3a0F2VnH3biBmHDGu1q/VHJPCz9B+T4UkVZevu1ArLhmcbr+6sdc
aGK5TI2qr+PTPn0yAkapsM0OEEFOMY0ahu7ZEALjFC5HN98+CQgu9xcYOg0aW8Uek7B9xqc/WR40
S+zS/b8fdTSk6xLgwlvkksQEam1PZ4cCFXqJQAqC614fMHBnpvXbNj7OKTYdoQ4FwGYbMnMV+0nA
uinTDCLtyOBi46ZjF+7e0wEkLaOKbqdLDOn0qiIJ620zdnGtfyYsidaWmKFiOhNf4nJMg2Da1eup
oSRVS1sNF1S/pl8qxEPnU/bmak2jrwi5L3PtqOWp7K/g8sn25VeMXOdrgSI3piVMWbnNk2QfQV6y
2AaV8Gook/GidWlkiSsF44wQ/eowTT2IeSctgB9JJrerjxDoG4gCkIJOPdT76q4AC8Z/S4ZZ06AJ
I3BB4RwwTCV0sToTuA4jTXsqgbQKFldV0b7b1bu3L4yark+syRAVci3pkYqCyCFCj6Cqg8428QnC
OGi42KEjg+geBRt8sbnu8N4CD3g0/mql1C3UY43mmbN6CP44PZluV4yjcTChC7oVhDoVOpie8xEu
a5XPUjLcw96p03l9S2/KAb/E2y+MOu8yzXraIptK9tELAtOHWPUaDohQUOqCudr9zrlxvdehxuia
JXSW00uV/eWeXlhDgV76/+ZPLpMqwNoNzVVLv3WCJ7R1z9a2ILAsqr74HI7hxw6eGQUeaUbysyli
oFnCQa81STZ/oOD3XqCoRCXWKNMdG0/H9w6Ld8qtrHdABNPxi87kTdXLdPN1pgRgHkKrQ5ofXY3L
DxsBZIWfw6dhaT3pWRahVvdDp7FHu7C+Rf3XHzWOZVlyxxKgzwSGGhDWcgAOK96xUFEC4nWGwwG1
kUu73/j5GttsZSyn9cQ/TWr0qbKbRs5tvD1OUVu3WS7eXJD9sieyZr2Qzxx7BjXurR5AyvSTtGpc
/z+leI5n21mQjMC3XzMpFKu/96azM1uP9C4sJ3vOLu4HzliuwLfJh+WXbAQ2CPtDxoUh3FmW+IG0
32D0a6HYKASl7s9/PUGU1zySCG3NwjjyZVrG+CvttUx2mfOCWA0IXJzZOMARStgmvBiEmtVRljlz
8G7WhWYY599aKgCF8ZfQy9B/y3jYTFcxl827Vdn41SgdRWtnVSQ7imD6vsYMp3bS6fFx29Thng2i
IhIN6wB6vEOa6QMyvVazGH229Z+aSige5snZ4S22vIUFdejr0COD/xAMIjKd08C9U2x6kYasphS4
UYFEGzLQyQuknr10tYEGI7kxQW0mBmZ5ftM6/g41gXkOkxgf1VVfuk7H6Ps7zGGav9O/lfUzYWOG
D3ZJoZWtC8Nbx7LOwVVg80J9LtxPF61NgwLfk7BF50IK8xq4K8jk4yrcDp4FrpL85sOgF21rj2CN
BijlvIHUksAjKGkiPjp+dpp9Y/lPectMTtsa+8oKrxOMIaKuQnZxHYMLxkCehybm4wWgAYBIaCGo
otUZLJMS1sOZtrYM4Kebz4WB3U2TS3tr8jzrvDzoR+I6VwqtJtkg7VFfRaKWBKN7mfXPua6tOfsg
6wJdbSU5fGzCCoGQ0VBE6qnYAhkfNbCRDT3hDnNJDUqV4C3fSVo5LC+OzvArrsT14XD9EWFAngi4
M1Pr39aquZ/ViNtFlp1JYJrhxJZAGSseRjPDdNFEkXOdI0wV9uNJNvzqrhl/dn4z5nIENzKn0ydj
72QTkiOaow0GN7OgJGfgD75GxweAVWPJISAE5oSDWYsSg8dnWBg51aZZJ5bE4RdyJbnI2HroSrvF
WPeNQqUbtutzD0bwHs1l67bs/osw94Xyskgr7p0aCrwlIflKAlBVPDQqNXfzMNxhqG2GZB6HsRhF
oauh0wxmzf1QBj8hjciuDDmfLVe10NPQ0733gXr+IS5QncG2Q/ow1FZzZJkNAf7DsUeB/fAfJEtE
bzLIA7HJNA15PdyRtdPMPdF+l1pYjHcjrcneMS3QdX5ck+MHFc3EMlhc1oE74R/91BwpvgD2ob1e
/Gjyll8BWiSF7B/Q2Nm6LaFzhoU39fx1OnOvZ6qbIm3kT9uXqpuonfOV/abGx+/mNdq4ITbtNzFd
gGmerNECCDfWd54C8nlEVdKE5IXRy+iuilooVKZ6dl4nhjrxzvaAPpuV3gLUfgrGKCuE2vFWHqnw
z5IHrhXG/gl4hNQZ/ysYNXXbEJSFf2eaCAL85wy8c1M85Bmq3eHRZp769kwqitJmN8c3JJGDnQUh
/3s5NliWaZfMt6mWfOpe0386tLWODtINk8YsD624yDsVrnASTZKPdI1J2JEN3Uy/FQAbSVB2l0ob
NYdu/cbzxvoEsNWFok4WGw/o7V9T5MEPtJEO+GxWBysCHhoyZDAYs0gbZOgnr38f9OeJiekiMhYG
BODzDWoR36qRO/2eiQph/7IDL/6wKb601Ghqzqiz2Mb2nqpj0Dk0Mj43bpdGheH2EfZzsh7G7hhE
JQPMo8QRO+OFMTIKllXUB4l2Qva4GwdzRMwgFFqNf2bMdKrUJJOOGe1HXBUEBtQNS2qiBjXedOrL
7IlBj8fEA2jS8/v8GdJY2ZBdkU59qqn1M7i1CXyz5lGARrkBHzc+9ivJUz/9wLFFLNeOE3Pft4Xa
/5fa7s+uOewjIU2t4na83eG8MPytImvMVag28KDESvCmcC/Dnk+WhWff+mDDZ6iV0MjD1eU6TkyZ
G45CGtZAgEYVfagdiSP6c9hI7HzAJXoojpFy0e2FVuWfTntiQ7qRehJtLfyIUrdvV97UNYivf0Xo
C+kLYlVP6KqZbUnWLWZNOqFQQFHH+BY25Dhm2EBhpGaFV9NE4q4ujFIgYI8I7PiNrQUOtp5pF3Ec
iTxELIvvYwteKAuTJaY73uyS86KPTzNh8t0IQt45C3Rp0ecy5RtVUhTNyeNWdlIVp1aVK5Gq6mtv
w49hGfVQcRwMxTJT24txvfRrCrVZUb5B1qLmdphxzZyVMqPqruHVn3r8VqjTWBNdHdzaf+Ylt7Fa
zZ+m0ia0fEkvWotR4/7KtZfLAKXAFWdIVRl3LyztM+L8+oJr+R0fvJ4Rxw096npO7U90cNcY3W5s
Z/m01vpjfUWSd8rKGlzgwYYzaAq6i06gy/NZKi/G/RCgwSbmvkyPliFkLacwECrNrlznQi8dIPSe
HGe2CoyKAWABqViGaPLvDL8J/rdThXGcKN4deFb3TkwbLWTueAlMIxDaVXy3K20P+i60EFeXfK9n
e3vKLZt1U4clLBH1Ndi6HgVH4LDK0BryPEa8uitPG0sw+Dl4nCDbYu9sQkmSCK2oFCnbq7Z+61MP
4dGlxFcIu7rDpu04J3ATG5ibn+x0W9+A/IQijIS2gaR1Ng7+vCNfzx+W309VSjAHZyNO7e6C1suL
zzWnqtiGeTiu2BCYORD4taiY788fUXYXvskyfNA3uKNoqadXoNY+JN7nCV88FpfAJu7MBN9GCajC
0yjGGt5T6itsRrb7ouMuf7Lq7D1d1geUOB64G02ZfMmFks/XY5B74bJzu8pk5Ktceygjz4FSZzRC
yenWp7Cpuws4pn12Oes4DZ0MAxryBlY8aqv+abCk8A3PqzPSd5erfbCmkSJCyYbQcXVLoRKXx7Dk
7ImeFFEyoE6V5oQYp6wmXqF/y8ThRLtxK+IC4vIyq9UkPSXUcAGg0oFt90epL9V1H3u+6If7Lvnd
XA4Vc/CuW3KnlHdqSvNcchKVFNxaH37gQfjTmkPGG3iadXtoEejlC69QDX+ooXDjKhJjyBLjVAre
H8S06/z6zvrb91avc4zW1/D3tNowh0yWdFKHBW+rVRPUAhtjtdkQX26o4q8pxKE2eP9FU0kB4Z+2
FUkgctWaTTC5aiHRae/MeHdQ/Y2UhtBrtkVRmv21X2IAEgciVBtN2DVzfX77dY8CyW6eNOjQY+fl
/cvXqM4ze+nUdDWUy/XZ2BE33CCRqlQcr4qWQReBQ53cvubz9XOz1lKq8YERHtWNdj0/QEqtuBMT
crov5/VoQLFypVEiTscp+B14VcJJRYTyCrAVcEC9u2ZytkJ1pY6yR+6ySj4WKxq2rHAg6s3t5f/8
wnJL/pd4K41W9S3bdkAzuQkGN7Tgtr++K2Hk38WOU7uGYpmR4N+YHHvHRM6vQlahMbLcqWKz6FBj
bg19gWcWbeVQ7juDmMVuQOR6qmpl3Qn5zOUVkyyBL180pLktYZjJIiZQcN9U0PUtOWbyZoP8cwob
57NKZOhZdHLP2khcPR4yRmd1Kwnb9iFN7OGKGroMNAPGDwEvm/n60gqugxijAidEW6m0zu1aeFk0
sVUD7SV7vte1SZzEwm1YsrCdHprb7LugrfLUP4hmJ7/+6stKAMBMU/7qAiG2v0TiTAycASaoEWxF
JRrSTuWIEypvoypcsx32hJUA1Y7wBYKyt1niBi3zozX6fVWXTingDKHbMBqoC3Ua76faESOf0SU0
z/hZNMkomsEOjAujIbZMNq9CvXojmU8XHBMIItYVUjJnJfi7HQxN+BwUVqa1xKOHV9DBI1UgU1Zh
RJWmjP6AceoaoPhQLokb8qpFtAirj+/iJmaPqdfu4QWRl4qJg68y40kf/LH7PM+7vDRKU4mHZuMV
6a+khd46VDuwih+H+F5PsOvqpuDitFmMi3tgFUEf7KZ1arRaYW2+i6ikQDFjk+OVIEYgN4TAyhbI
kZ31Sbf7vBtSSBMTn7igM7CIlpyc6UtXez6ifqXLRjoMdItGb88c2lVbj/sspgKFzmcDrR37bW9f
zPryQAHDT3kKqCSZD2va/KU1PmYhhNz9KYD7vQCntveg4d8Zc/VQn3VQZWhwTx+rsnsM7hM5ILwa
JhS75i74KqhXUbY17W9Uh2gulDAJpJJWrX69gvS9DfXUqpzl+Jytoe6k6XePpZQaeAQWM97srv2v
YXdzBUybNUMdgDtWGP6c1PrzPTGDKdMXi/GDi10u7WvZ9l76lZG1uCwQ40Oqa80UbEq0Teif3OaS
O0pQhT++6nmUHPZCjfAxz6a7Fl8qBQxNqtWOh1MEJzo5m6Foi8WAzhhc0TB7/TFfdrJOPnlypzor
9odzekKbyVCc+Iy+zCKokNz6YXoXEQcre8sHiLjCE7jPmD9Yn6mj0v4ASCHmHKQ1UXfevhmSYcep
B1I+RxZ8bUIMVo1LtW5X18IDEv3h8eG8i/1/8bfyCjKVqfo3vTuiYKBil6jzxke03AmkRj5LDOn5
nNp7j9na1tPB5Uz+QVXY7ZnDixlk9NxfjeBCyHW81LnK/x2TEuzUxZWKGyvChLBJRC5S4YZ4E0Ss
XokpqiVJsn4aP24D/LAi1lUrpp/mRL4+LTux9oCcIsodmbodeuUh02Dn8YakIHMPJXhNH8YPy/CF
DartC+OSruLUKA0W2o67aMPePdCqTJzJyuQbkPrSuJaHAX6nvEVHFsWXAPJwWdYz111sX6o7qv3w
bom8bobGgFwBoiZbAB/XFCVQKXo/p5tybfXoRHXB1DSH6cxCLrcmPn24xD0fHzeVx0Qp6Rt0iIDd
XAHgiuujG8M3dssTm/pw10eLflFbO8uFxnU/jXTATEmi14J80Q35UzjpTlDkr2BxzTH1y6r5Wumb
NOnzchMVKEY4JhpZ84zyFgEmjYYjKdTJgECLcRh+gSnB1XH0reqQUzLV12PtPWxuJcSvzMZuHu+b
jO2FiXCrrrFbK5riRL1Mm+QCw1tvNDzeNvyiUaA9FzXq9qttsfSHOFwCq614bK+QVlV6PHvT/xFZ
SZdTbDiD9m9u/BJfdXoboM1Bs7yKG1W+VXBOxlZbaohmh41F8YfKyi7JBMwhuGP8XSyc3iRnPSNl
2SwrCRqHEhSDI5fBNVVFKOJnzH55+aECGhAHzUva5rIRXHWnV+nxtMceSKYy7m3qJUy+DCJTuDv6
bXuOEXdYm8AAH43lHjHUXMT//2rQmfEnm8ACEHMRgIdrRHcO+g2/ww2/EK6q8wMivXN8P1FNcgsf
W4V1zoWspys6+V1HeONiSNgjV8/qIDPghOyy8n4fms6e9DjdN3+qdp1vnEAfNZx4ttfNjMsxpeSH
mbB7OTZ4NfyTAH1MROfhFGrpuLAVcsTsGuGuxpMsCiZzl3La3h36Fk/412ioUn9sg7uLKmddqBfC
C8AkNTxkqCA3YV8yNHpawSGdJOPJd5pj+AI9SxnggUG5AGxUSabs+gp24O0kapHLS0jIz3xL5XMl
s5rd3LaTcIV4E2DiB687Bl9UvEJgezR9pxw8MXsoo3KKyw5D173y9DtViZXL0mFnJm8X+aSr6qGh
rW99xR+oH1h4Vrwey6ws1HbGntlGdd+N7+M/SiLVeI/q2yu819UMXr/RK+yMWPQklJR/9NtmO/XY
BNvQmwOL2T4YBXu5t3BHtrnTbEHEAWNQpqP9fXjwDKrFXvJBHdhNN/7c9bhNtZGSQD/tA3fXSqdK
DxMLZ8SgsLFsTaNQghhC5Wpz17G7TdLN1Fgjkr1zLgZ2POrgubm7CMpmDV2DUnOA/1JgbVD7ixJm
D1xUQjEi4yZAhobYuwWQ9Wg5Y7No7jR3jiN20UAfVSxG9VwWQUJUP69KieM9ucLrNeq+9T41YTDR
KRaL+fL1Vik/9EbE+HbVqsBH+ygRiXX0kRSHFe5wE9nbdMbH1sZghlB4UWn4pmrmF260NDo694Ny
ewyHywayW0x789zFvp5FAay8s45Y2/dZH0lfTBzjGCdwZKxTvdstOZqtVhY6iRbJoSlC6ZEkOfj9
ah/RsnguprDFVGoYJd6VYJkYs3caL7sHHaAeKcpXqCnOYuIqChKFJFfYtLemWaE7GeVZbRh+kN79
w/pwF3kYkenVveus6FzKngsf3xNS+FOuY9pvwdEMgpwJ9OBqF7SxxqtQJu8ErRepeAzE5mS15HyU
tVNsL5sqf9wW8bG2N/ov7bm3rTyIyanbTb22g8GDx/rFIGxm6iljMMHWWu/id3KClzwyIzWThLmi
2UF7388I0hvYatE5Df5wUPBby2tGRlIU3B1cM7hwl2prt0AiZZ1FdJr0oAoSFUzzbhS8Thv9dqqV
uJFBk9F9wulOyeMgIN8JiFsiTFeCoAOgShxIkM+M3QL6tCWn4Dm9LgApLEuH7piAK/sGBhHdffJv
jrkCXJtE0gtaAraWFMpd8ruOhf7DSjTbQRJG2NZogcEII8F4JLdQhn7ha0ihKkwZoJs4At2KWAZR
HQIKq2b5XRxSgls2nehbCKiZCo8AmY12D+BjurAPnX7eBiO2YNRZnbWb3ddLo5l6tgqUG8XAoRiL
Tse/DbPma9kIPjwiX2I5cMjlrZ/RtWpDT4XqCauOh4IQ4w9ve+8fWVDLMlZJSy7nIpdq8fo1uLIi
PvOb5brj7Tkru7Mj0/XV5BkTpAvw5rK3VJEqARXJrqQeYIirHpwJLDt+oz72vOTY0KVRt2SfmYEU
yorksK9hVZ24vQY+3QN3rV+yGlxbFDVDvNf6hnAPg2BlgileCZzz7mh0PmNmUqCh973L0DdyeDRH
wRBwdBp1wzSfNsHqpyRSD7Iriglxtv2wSfUorwe1iKJlXJaDVV914lIhgOG/qqHX/2VLdR+xv4/C
3G9cs6PDLSzwdwxRz4G1jeDL8/CBRuMvevXAniIqkKxyMbPKPw+ivmmKhHAx58QpWaUxEYvIY4bM
lEJhtiYsfr09uC3Qy0lUnz6iooBhHO0sGOpya9OJLkZqXzw451PP1xzsiAWeN7YB+By8YJOh0S8K
llaNQHYTZF0dMeTEtySAuqa6ZLbMkrBWt3Rh7hQL9OrI0CKNKYWcIxA8JDhLMSPLGQmuXr93ZWKM
Z7n2QpuOwpKGYV23Rh6UXIgJLYGrfxhKw6QCwTASoJb0OJRL8tg527RF7hxOlwg2tcmXd6x0Wnw8
aObDAC3dWJ6WuSwQBz7z593G+7Izg0VdUOhNmpW7aHkaJXY4lzrnWGGMyCtjfhLceOIo3IbU1sZh
3Qoc3Eg2jfLK8cI/xIpvkzUge6iCnsbLIT5iOH2p3LKHQ9qKFPTpcIoTj5YZSpKXkjD9lYmWlgh+
IPigYXg561AjPGbBdn0+tS4+MqEKfTQmNYAtB7r1/EtB+km5pog8LVAPsAkkLsRrfnjfEOunUYnd
U3Vo9JozC5jQtUG7GNanN1eBXPIlEOgSPmjcjW/M9tCcgV/Ysn6CeKlcHNEh7YW4SwTKi/4d4Baz
eadswxCdQ6T1G9DgInUTurOHaQtEVsEoxRMxQAhKxv1rSwhkk9Tm/hHShipDVtkCtReDYeIYhyPa
JDBPW2OcarRgtZs9ckxHt0JWK/D82fLHM0CkEYRm/QPIQupB5692PuVIqXnPqL8uMO7hS8m+qHPN
df+b/kep6AHppSe9phXXF3P4UT9p3JgdAxBHzHSAcm4FUuseEXryqkAVS2IdMxVTNWxgjbOIQ5M9
b3J0hYn4zNd0y9jpBdEqHl3J45djpM+MRct+yi2onYaq4mCvi+AO7IJuFA9Mp785eU0k511nb1vb
xGZisMzaujZjaacDkhH8uMUKl4cqJz/VwVxKAXoD8Xucwjhuq2+/+gSbGIkhRF86uND3LZv6jJc3
NjJa51++sOv56ZScSEgPT2VKDT5XbnAFTjCobWm0L6KSyAQxZmGGmjCJyDJDAgQI8o/HAojDl/S3
+TkM1DtyOsIp44GHPL35GExLipNANY++vGCqgUfHOYqr4kEtdfTjPtJD9PDY3EcLoEkW4ys90YPo
Q7Nv0gREUmAEJZa3+JteYvKLEcU69K7MCYn7k0lZ2MtP0/NnQ8Go6EooTCYEEOqJYReeHCqtUlQS
pcxuzD65BpduWzwdq7ThQjYxjC/KJv9d/A8jkQnD1scJ5hr6WLk9OyzPspSrWLiNCRLn31OhEOKj
gMj+oEptpTvKXNoQoS+RCec82CaTKOmIZ7FEi5PI2w4Rzo3oeWpof/8gWgXT1zQKHP0zd2w60l5X
sw2CyEUcfOyysY/NwTUk4Qe4K0Y4uQIIyLCT0GmFIvLx9hgoENtqFV8GV1qc2b+3hRodjn138775
7sk7fA2dfz/DcfiCFTHbGxa0w/LQiXwD2fqpddsMEeWyU+MjrsZxkxTbKdEDSPGrGEqPfF5JqYOI
LBEQ6jMOtPPSnLQj/mQ+AQWHiNKgLG4XhvZPonxpOoxlaDClrys2PYyDHf82jinJKPRGfWL86SOC
mYswpLLz/5NgT/a4GdvN0aq/NXIpWNt88QVrjZrbaIhhTNMyj2hJf1ngF6+OrKTUXCMkAgaLgBbf
WpunPy43yaIUXi/9zUJvW+ZiGr8Qn+Fwp90K259VxlyoMoDAZIJXXK76kdfq/PWGKSiQvEzFcqxT
iu7Z8Vzp2D/Xu+PB6KLkCDkFES3l2bV0qGfIH1nX/S/QzMQn1VnXNpXTjbJOovdggRCPqeDNrD2z
qJJxtjCJ+miO/BObXKY2NcOCdVwH0s6mcn0k5JGpdRTwEkJjirSaYTsAnk0nPKbt+F9sBpcWcmxG
Me/7tK3CRql/jyfdlMWLZCOi/5coAMRY2GMyQ15zFbYxPXeCXI0QWiQH9pQT5RxZpPcjLfcllmXJ
7UDafbIBKX+dxE1Sy7qd72h8zwgQo7n1LGyfJ9RMz7tpDMhGC41qKNXEsFJyCN8MdtaWx+/qfCRx
pc7q4LPnhplyNYgfjlETXMVpgmDRoOeadEjJQAcIXZztO1LQJ56g4ksGPn7NXdDCs1hf2qCY7AKM
mUX+x/2mLUWHzZBFXf5MDoA6ffJ+otaf2IDTvAaMJwNQ/HthtjXPhlIGi5RcFFLlsJ+z6zXBWB6O
Qi1nhyMMMEsAfxUrrZKAG+feSUZwOJ1ILfE8Vu2/NpZuMGU6LvHokIwg9iAc1DG6gswbOxv9lT7+
IzefGLrehEspfIKqL09keqGmaEjuKk65iYmiNSkSieyM1mWKdRmVd+v36RZForPmTPAw/eeccznj
vI3SF5/jYxmCblUKdEvsmgTNHPGck4gd5Loj8MfckE37jel92JbNNHmHMdWdB22NSO3XUDHrebp/
dL9rkJJ9YqfpJL4ALnd6jwODsmu7EgupoNU7hvTZ4+ptFyMkjmS3ec9w+IeoHaWoMqA1lN8mowx4
ecnVgNbsae9qgN9zONvykdL1kunXiKxr5m248SYitLMg8VZkLXn2eVBPeUlUWfYMb1u4qXT1/tih
h+PsSeQAEw+eB9ahHngARTotd59IZeTnlQSKvYc5NChpTY32H7dOAXn2BYPLb8ibQjWlRX1/mMSM
kjGxTE3QzHBMoQgVZgXfmy4Gku3OGBvFCYxtyPs27IzqxMb41LCPGr71ZNGlXWiwC58ArG5TNSaG
PkwwEvL4i1VQ0TQsCb3k6FsCN0dEPmKpxZ2GcJYmW9PkvJT5Vm6Fsj6o3GfcHw26TaXpfpiRex+8
Kv0w0fnhq9ZdRbH7G5vd5CsbZTi2mafe+nvD5KZCYHtojIKevuhHFLB3HXOph0lgGoWl6KEEjHaI
tWZ5ef13dSfu1JDGDOhjtxikWTBl71VaKBmXS+4xrH/2fgpkkn7fvkJHsANGvsImiwEpxCyGNdjy
yizIWrgCONh8r51QmTCatLI8fulv1x2xpmWb4pKwYrPClz+8TPcIoKBTAu7aFp9UiJEUsskHLFwI
J3ih0wrjVQ2ZwzoHt19+pJ5Rvl0OUe4ZviRduSBZ/s/bDjSvnb9E7h38sD2+GHYxn6Zv5MJM99M7
y9rPC7fUvUY0oLmKBGHx86OPJ8tMfH3p2vIfLMTD7XJW+Vk8BnuHxmLvFyV2yhSs2prr1/uItOwc
0Tr80+laeYyy7s+QN8J0gigePhRjAgVpP4qiwOKa3WlRDqSkL7Ayi9zE0fdcMRA6X0yhDQtMRb78
saIvnvkt9qa6BALT6R9O+h+qyQ97Dg62c7MyDZFuR0LK4z87NFN4ybqu8wF464BWO7Vf22GcdifN
A0CCG93aMG/DkgBYUPVKL3+68IUF3cJ9yGLGM+yGjUV4T3fmqjOWBLKzIzI1CRmBGEpixiaWfDGe
7ucOak9ulfd0f5mnP5DYa1zLMNo1wVcwO34v8CFs+0Nnttmm1SIMWpIGO/6XGGLgRRKFWArr4+hz
OCqwqvAjtBev8CgYSFnU5gp80Td5VoWnvHRYXlhPVyAy8T4LDANSNLDPhjuYYRtgaFNuCZbnMt+G
+DssQ+LXLT/MEo9IH/k5KWJZsVB0peYX59eKOwx1hAlfVThjIlmz0Y457OtRLrjnY7I3ZUwmWiOW
O2XfmknC3Yjm4RK/i9thLd5T21kEJlqOr1ulmST1KJTXPhfx7doxC5pjPrWQikHQMeE1P2Ca013L
GT2gENIZtFU4NGQW7KNWRCZaTS91CLEIXpZxVsC8LZw30Gy9DimO4GiZeLibZt1vcwXfkJ8eIDm1
i5Ae66QJoPJqUKr6YaNucGYyt4xTAwTMQ94gZkWEy9et1fkc77Ihq7hLEUfdVq0x1ZHgtkq/PLaJ
nvQ9qMd48fFe96SmGoBrGFKSEVwViy3pGrtdSLvmklcYqnIKKOgqa0/GBVMKKGFDacgeEqhJ+nJA
mSz+kK8D5Wh+WxH56bw2qGQkUIuMGP7o54P+DMuD5Euz9/YLpgt7oIVFAFRMEGWLIjHyJBeaYgm9
HxYG1Cycq3BmA+BQusATa/w5ZDVeLXrvKmZlS7waaAdRPBJ1i20vlycjmTNpfNyRf9FbuHdFoAvF
+hz81y391vQobJ+kj2TVcK41TIoV0gqLXSTRUlqI9aNatwSQJpVKVVQhF+kpzKP4Tb2kx/nYiYUD
JENf6jk1hbISbZPQ/+9CIzkuXxCDxgMPjD6oS1L9v7c5vXzPgH9PosImZ4jCYPUNTYokngkOBbGN
9zkmrUtnQZQEuhVFul2Z20dadx8a1G7be9Uf+1n6MtnOISOuJtZZFL66Vjr96WDEmTn0kneEhzeA
MZmkVkpBCnyVu2XGKs6D31WS0TZv2VNMXVs/zs2l8L1wRYSnBllrNqiUdcaRx62ZcuzO6WHbh1oh
pbjxrttbeAzECJhCJFbsH+ECBN+HcHfT3BJ8clNt914cF5CqiDEtChBhfAxI+0ZGKpNVe2ywSjYo
VgZ/+CsxQL7A3q1gvnkGkdB3SAwIUV2lfZanVUzVdbxDJx/z/NFHYaP2PhlYjKaA0AxyEZmEttVs
sIOSY5WW86/bqwMm8myO6CGJpkSKvbC0BuAPSxr/syrM7JwO7dXNZk8xNtHOY3JfigJxijB8En1J
ejeziJIuQe2hLwVekuxCPz15nEBVLxJzf3DEARqqxbwJhMZ+xuc3uoWmropwHXgUT+8cSYzlezIv
0/cvqIkbf+qFPYVYaTvPWIjRUeV3f321hYaXp0GS9K6dW2XSA6WNWhzdoyCypr3N2g06m6OEr06R
62mplEv2k96Zfo2QrHW5UJIsg1UK4O+4DhBqfAqvevjhK5JBypyTvTNkdL6q4AbqSzuASXVEbfG6
V5luSGrRcSxVZUzzXKY3jhDxOxjcfLJ7RWpHbfw1bK1ggq7yBl1uQyQSXDGe7vId1j0dMxoBDLyH
qfMuCaAnFz1pHaICJQ59HDDw72jrS6GEpQESej0O/TsSVLwngAwk3SBnV8JvehilpWtkgHgIzzrI
6OBp/H7V4dXx1hIXT8Rh9dRdrZtCrduiCPa+kn43eUDWkky30oaSmbuHDvhes34kMp6Dowfnx74Y
6eGqPSyzpnXF/H9AY6PQZCJntvbXpa0a9I7UEyfXR6B7jmdYAZsXnG4DIhDQZDe81JbKDVT+15zu
/9NGwyrSuiUjVvKE5lnD3ee6w/rfdgkOwyDC/ifSLGH+U9nd9utRFvm/UA0sAGQ14S29W1QHxYj/
5trJfFFYNQqk8b/IaqWY2A5uB1g7McYyUxDhe9RNIguMJjHuianmBphGkJHlwc7d9lKSSPY4N71X
ikCFTaQi7uyAhR+qcxt28pazjojLk7I/68lAx4gaAxaJmfX0iLWjfXQ2ZKFsa8a6yjODpjN4ENeR
li6lEWzf01b7NrSJWZYDDC8G0tf+o+BbuVsBGu7dk3D87sBMubdPBNei4X1vL2/PZevHM5s+LV1s
mUFy2INeQtYMosCfE79erCP9QNAigsFUuc/laI/q9rgnHvsCoR7zUbBIk+t4ExOYKhDPPnV5v0Kd
7H9ymMv2YoIO2tnL8dKwwyzeAErWHZ/5QFP4g4jCkyXDSV0va7W+ouytrhIfUQYXvOl74irMMmUs
qAc3QucZwCRVmjqP/GIQnz0G2ibRxEWTUishULvHbfSnokO4JZMGryYol5Abt/PD+6jXeTUauuZh
FnQ3QPkxhjzY0ONl5K9lEjhciiHwIqpOPiQfRR4j5UK1N93Iqo8J5G50LSIOVXSsOiSyMp9Jc2tU
iWzYzID3FHKEM4p1MKLQyCgj3u4giWNxvFTzyY3dhqS0rBYv+WBNc9WTMkL8q3Hy1Km0xzNmQy60
EutrV+1PLgVSma7aSsczdZkSYlWSLgeZcFqmOih4vZ1tWmD3MkUCrYKd0PcCV8IUkgQIxR0og0zL
Xv5+eLoene218HKi+eaVM6jmCbendbpAltrUldKMXqnlU3+DqVbaOjrUBjLsHJ3JVHeDfcF7PPW5
02ZdgH/I0Mf9M6/dLRryWDCZhPny91DGlV3F0lIGrrTEI/kqUczHZJFDrQqbsBzNXUH902lwynCT
CLypNs0g3BDDAmDvmiGomUdc5ySiBpsbPgAPlcr3pXCgbcdYIDzU3F1dKsyQPyUx2LBKA4t8MU0j
reFxwrPXdKQEo1AjjXCIG9CCkjf1PUA2aZxXzB3DQ+YkTXLWFJATRF6jS1pg768OG3S2/2hIb07B
Y1iN9Vrui9DMQiMURMeAUSN9078Nw9vxg8rbhadw2wdLcpe+bdXnfM+P4/UlU8FZM0vccckOZm5t
KmP8bs6wBH8BPCG/gNxQ5/eKsjc7dWhRzXlRo9K9hqstR6FgCmIIaNBmZ39oX2u2NRqanUDAXJXK
D25xxUpcEW+MpyJDsRgIYXkmRMVbP/XoR1/o70LY/rnhALfMa6BX1TsyEn9MCAv1suzo6+cCeuUT
7rkiQ8wsTWbIokqvADt7n6A1F17HjYAKqUmjtuUOjqgiz6E1DxH9rY+b5MUJ1S21HhRf2Am8ukC+
ELCw7EPu9ugCyeOwPTrf5eMwG2b9JT8wmGOy7lmb6jHnL/f2FkExmRLT9sVsHiYUS4ERgCmW3Esm
ha0LRExDvR9/pkZG3oklaRO5igh7ImbymvSWN19C0XlMvryWDP5tivssKeVJ1rIPYcMzLlF3ipzc
ruvXmJBDZnzvVLt0zvDYvsw5dD7IFsaktG6gzfOIDnCqr+4r7vAzbjQVGJ20EJPIuEbQncNgBuIz
rXc4Ca0uw9ixeRzYkG29F3ytWE+JYUyrnQW+LOrokkFM+wrt0fJyeurBwmFNT7lMBp3ET1obm0mV
yWHCDtfmGMBXASZOZv+5Yavf2W8xfQobxwlHoQ9E1Yw823023M2V35b8ueBVHg1sj2wozJfPh0d5
klTI4s42TFMIkFmY2fxjAqM/SbZVFPVZnzhCdY4bllK9OxD8jnvjtINrjhCnN/mhoX3G9ZGTRsbF
uqzzixOgSdxp/63i+74dOl8cv67kSC4RBEARE8AnRu6aEP8TwRSik/l4PCWJ5qs0zjL1c6TdrqEP
zAuMpDNJQHwZHDph9zq9PG1luAWDYOtg0yMK3vFAeNS8uk9glrLfNPvBSSgV/Wr9A6L+apB8TK7i
EzmOluC9VjHdkU8PXEGnFeRbTa+B4eSM4xKj0Wv9Kzju6DQ4F5rXDGPZMv4iXDDhuMYT0fOMLw86
s62RXBG/FC8BfTg5ftKs0Ker/06VcF9ElX9x+QfDEmnefWlK8m3CUv1C5VibBdI4d0hA5I7JGwOm
ylZZyuLFn98kW54xlE1j8T3NhRvYqeCEmDgiN/lDj7BBbJJvaJvKDMUTVcmUhdeLFuywgLHOrCfG
ApOyfYgvzin2UdKCBeAgz19RpGbFCFzgLCsSVQYU25QA/aRDL4a4Mp4lovIQSUo2e3AZl8iSOduJ
o6e5qI7CgelS6GuqDgn+/3+TwFzbMz4Y8UBij2TkwLvOInW+Qy0kvCosNzhip4JUqCH+ObNk7LJt
/VfoE8eS622KBEy/Pgu0Owi7FThMfAnfrIn5z2dwx/Eur9/V04PyiEj4evngRyOe98kJken26Oo2
l5Ot9RdZTJIqU4KRVaLcgkVc8g68eNQ700uHPF+3x20Sw0cjHpOn2qPPsl65mqL359I0qwCZjzV1
SL0UQVeYX4+/kx8CjWsHxBWLrAEWwQePxlNEXCh7WqFNwAwMjEzXQay3N16VYGpMKD/m9nlzmSK8
cZXvKfwkS+PnWXOIoJ3kcOdYZMQuyWilB8gtR1v9dTYtozI23EuwgIAqe3sI8/JJeM8frXm2ImJ7
92w6ii3QogCamj70QQbMnaoasL0U0sMZbgtMSkdlpLuVktwcYripYmNphFljPvCXgp3TOuALqxJR
svsYXztWrhM+iQcg17E2IxgAEuZP7tf787hmBglndJpp9f59RGI+/ycGZlyAMJPchPdDn1s3ZYYh
123uJXjq3N5FuZw7VBa9jhzY/xynBypOaeXbs2sXEV3B2YffSJsdDE83nmb2WIegDaDg+0Szyta/
0YbutJq5Yv3ztqxZsbp1mxe0MSGW3gHc0UwwwgQnCpxlm0BhhV/q+/wE1q8Up5HPTZy0ulafqAhm
GoEMgdWJWU3u649hEwpusfKA/Bx3PqtEvyq5LHkc/4Vy1OjxVwJA9AZmUEtnfBkpK2HyzkzOUfaY
c9cojtbFmiq9RInVMck5PybLvNRAjpcoTR9pnXT/YzqdqZvhsD3CmMS93QxRtcNcTO1sYqFDWdKE
KH5YjLBYu0Q/utwavFE4gOgeZeQCjp8I61mLGtHmgxC4LRmKDPfu0DEWtqXLlje0aIcNP8fxKLvj
pRQlNEq1lSHvEvlFsQejRkU2nm8pxn1zTt1VQ0cFwhMYOIj0yO2bdvFaq5VDRxK7RNvAXmLomU/J
tX1mJqInZ0MakOeT/TC+5XlfxIR8b33EcgcOBD5IU7SCg9eQp/imCMqexw6RMLHCWghsw3igK3zz
iSLKjAd6c7ieEO0Uz1yge6CWS/jy5y9mhAVDKF7DleMdpBQJ11dwHlgZh0vY90SMFPB5ahJB56AU
CW06zSussCac1v6F7K2Vh+wMsqmU7jSFl5AjxHI82HuOEqUOFCTGBELcxXAPm1DNPOrqb/VC1sBU
3EJ41cPWKXRgTI3mPFb3TekvnnTn4jS29/IOCjlRUbr9edDsVcUT9jmj+OS/zsYCX96P+GFMObK5
e8ey22Ja0NSg0gCngHtzLRn2fssRHkPMCpl9mcJQhyM/vhJwUn5patPT9m/143qpdyTDsVjFy5Yk
GUkjGLkL8+QYZR9I68zUqnuBwtvPvRbgMdr6ZknHnw75r/2yetMrEfoFPMEKE2ot375/qJ6WUQxp
E+EhAj/TRGD4qjyNoeyXj8mCweLuql2W0CUTWrQYEa4/hSUNcXUnLl5O95T5poGf9HDHurr7Gx5p
lMFaYqXXo+Lo1KYTDoLy3pmQt6sqjyGe4uzincf1uiCrA3aJr/UiFwAP174HwZejol9WchPkP8Jb
Q4KwImEuz0UZe05jBUupx6nUH0tdml9CX1svs2Za1xdLs/j6OUY2oLAd/MeLE3qNSZuC7r/cbog1
ScI04ZiAI74eK//rqa49XXVtm8I0OJnETIV5UvfIwVU6BYmfOOTtixlJjD+CW7UpxO3UMjeOVv3b
Rz/VtUaoqzDe1WVk/DqXaJBIZ6d6qO7TdPYhaU7YhU6D0EvFH4wnLC7lXDw3U1tTcFWJ/Qv4rnOV
PJNJHewXrOxT2o290oQTqaZz6XI/Yyjs8v8A6IX0id/sUbf9rU8l6FXyUCqwnlsiX0lbyWI/CY98
L0BTrNNU3Yjdzaf6MHPs5X658qbxB5ndH2tCddu99klH+ohU92d0VuLoxdR/vPGIjSpT0bVedQ0U
xOrjj8B0IGQpkHk7hcHzPtOD+QtcHs9oAZkQiaeBRGFpYHr82m32Txht0E+bIPDEInbi85EaQaDq
/lMH7fzyHLYhzAACpvIfDLe5uZACDUCJL1uY2GxQo5ADxlu5rSz8+gxjtJXv63uPPKBfRTmxorxJ
JSthu60Bh9gY1xL4gx2ZaeHhAt8M3Gvx5kCbYfGAyZJ0oS7NBnCiiFwI8EQTrK63j8aJbha0pCy1
4Flb9Ri6hxF2D3fef01FsdFwGUhMPC8zM24CyCepbiix3kXF3HXiPpe1pZ3xliUC+3JoLFCqUYd4
1/xTtbDLxEg7vgzcgzOKv6o1U82R2qq2Ypxg7IIA2Gv+zTAx3fR8xdBE3dUzjbZLc2CI02nXZJcO
pTC2HlBGOLeCm16zpwuRV2MngnNLXwfwrbmlf5atekEnkammCPbwvMNhvlZj+VsTvcGQ3NA1oG6d
XqjFlAq1wE9MwIHkEtDyY5LGVggc/uzqMhRbdJjIyuwYWikG7LIJEkwXj1a0dLXBnQM3ewg1oKU9
ETxCd5VpXNymXExP9jNzpze/EbSXbBNommfRhMBnthW9aBKF/pEe4H+bRIh8aJut3s/f/kpji0LO
PaDHASfi+2AvSL0BmWFZlYzmYAThNoAy+SrlKB24dTmGnsmNWEnQJQM/L+j9Qp47T42HOESU2g8o
yLj8AsGjpjTDMTEkysqiZp+CpLvNYlD/DeCnqF7hOesAdJ44Jy76e3OeE+737S+qlefW/yP/ZQwv
QJ5t1De5TSN0in1BTNtQmv371N5TYATbUFt/+B7uXp+A6xCzzywjwLHzBDQ26mftq3D+az6JGOu2
BDPstyOVgDeTraGcWVut66h8fyIojxcDGGarIzeJWah23jUo1K6glGh7zEoYSCdOtHd0Ngw/AB/y
AsrL0CGwrw3rw7TfM60be9Iw1r3r02JSHWvYK5wCQe/NmUYtaaw4uWMiGudNkFv1ryKj1HBXnOZF
preICvRJ6tMgwbkWPjYrmVXTv6JgUjby4+vMJxkJyiRVZU+O+xFbyVKKKMbnNvZfLIJGJWB8b49c
RA47t0Fg7SCfuvTXfsDgSkBuvegNcijsa9QA7al8GJ9MWTb5bt/ddxaRCpXoXpdInJnox4Zd8stD
1s/vvsuLGn8gXG3MqUar4Sn0bVWRFm4A3OTt5xAED1PX4OfrukR/wSSD3YxTbNEJv4yGFIAfz8kR
9KM6AxYaVQTwrYmQJ46Sn2RgtilXGph5Of1TNOvbnSr63OIX5M89dqslUqO92LXVJ7b3B+0B4QAZ
FrqOeTllYDEA10jvoZRUr938gy1/7/lkzn4Ea7MpTv8uxz3pOScDTCz82rT6s0DvOCuXQVi+wU6Q
SMPKpj+RbEXO2Jj9Fr9rcm9c76v+CIlju+REVsJpaCxOeTYO0sOffBYYvjuA5QHNm96HoOgUKSvW
/Z8K//DEVyqm9OLyxUQyGv8wUMIaFP8Q9h6PnqqRTZ6X6w71HARyel4yZB/hxDsEb4g/iLRSZHyb
3LkMBWe9EzMmirTmM5yf+yGRixmc1xFfRnUsaZqhGYCUXvxqTWarc2yS/6+8762igjVxRTHwVSui
p05eZIV02oBvPTjmFessJkil0xMqpqsy9YT8nkmq9Q15a7R5iUI0p4Jnm3lzDZ/VgznK1lUqoQgW
N+hWnvJ1gDk28xe4xLcGNs2OMDS02/OfbJaTFY4bm+zaWLcXCDc9eimkafwEt6X+YJDZM7QzXxVs
DcSPd6Jy0kv/tO8Dm3e9jaSXuS7WQ2YDQ6oBXfQBAahFj5WqsSTnJrypsawe9Mf0G/NTG8F6TsmT
M8D6xqle19MFo0NIQX2lII90ZO3Z9ZPG70z5pTB98GsGcEXH7ZgT5VXXHIITrZCsqpoivMOH4/D6
7ljWdkZTJmbLh1OA73uzu/DokfAp3YA5Gg7tnvfzoykereHq9RB22NdxyaLfDaostN4rh3mExB3g
xCRbvlr6p0iME0LmGUnEpNkAz+4R5siKtZRWGSEOG97JEyiNXUTI6QbZrKG04glORdRW4H6A9pxm
GBJwK81YcL7gO4sGy2mH4sntbyc25j6GykGHqCoKz2KWH+TYSERdK547glbKKGGbcG9igoLNKgp3
Zu6olY5l8tnFZUibxmTWO4eZ2lgdozGPKK+2g9UCPhiFzVR13VdHhK21i1X+ryw7lK32Y3mtINK0
UxvzbVMnqUovoqER5Qeg/nh7EMsqwrOovrjIap2ry3166FPPqJnsGddkHnMYzeREqp+C1juYXYZD
JZKTJV6hqQanx3FQUCicHueikUXy2q9+bxQXyS3QBibOgD8wuT7AR21+um9dTRMwke7Lm3MHY7sx
3kzf5uMKwA6pi8eyreCS5Z5JhFUO0pMZLmKN/qh9feuFv3zeXwkF3M4VwOZrQPnpoxUEMWSmPGCn
4tys4MQOy3Ye8rMSUiWY06A1eGbrFOuUd49VNNLMhstLIJEojt5GO8MfLRD2EgGmgju7v4D2SesI
SIVXnYWdUjfbOY3X9EpxkGuNzxXezEVo1ZnfGviKcz7+/GMnvu18mZDzaImq8F4fkM9kiycp0QRM
zz+lwOKXmhqnk1D3bZ/Xs9zL89h0wQdYz3elXaZ8TYiHqR3ZdYUYcIDE2JfyentO9igOyTZ7D8B2
RvfRj052v2sHLd0lbBqLqgKpr9f3vzyjK8KgEF4rDaTsU4eHOgacCVpzeKgAXgkZO/rmH7SHiBPj
1KVfm3tQSFWcyt7OPlIxnXKzdGGFC53hBssNcKV8fIGkI3big9s0OnvorfqloQosrNRDxfDzMCWE
w7ed0Bxk3N3/AXPLB0uxaF7s3+AS2fJtrY0G9+G0S9nwljMurijyobbpMBXagRGNJJMmIFzYDrYL
dTGT5muKSfiOPgWTsGYAWvXlBppKEEjl2592EBQ+1P8+YIv5P1yKlPQzNYQued8gssWon9RrFP4S
LIuraFdZMwosVQFYyVfWIo9uW3l/VyRnYgmu4AWbihBS6T8GBR6AFJ5tJx/pnPhgwi42KwNclJOo
dwG0EHTDiOpA8tgK/PXYvlHEqyATm495T04F2qmLnzwl0xU9z2t0kWl2hRvacbDozX8qoNqTo3jh
6SM7vwZRIl+4dM6nrOYuxN+TGfGvjjPOR+t3DiKlKUQSECEUTVLwvMT57KtBuq4l8KTgO0fUEXDD
pUjWxlLyLf2587JKbQ3BOOKnN7OI8D6LDYUWDhvSIRhcxVs1/5gMM2Hu10tg6CWpSwW/Fyljd1MV
MhbLsdVTXAzIEmxNTLlNcTxzPTpd/vsyJ0r94YBFNA8qWSbVblpGSPruJ5YSMNP0Xl0imxBrlwCn
03UQ6jT9OiXNibVObsGZjOBXEeoOYrxA7tgcd4BnlVLZryia+5afplrzBu2MwC2GP1D/rGByhkm0
Rvj1SeE1Nzn/lz2wcXV9qthn5P03IDAeduLec6kIXo8DG4mQNbrlg8N8CTyXaCN6cYQRI0k60e2j
jaoOYrTEI62+bOXClXnyG+wvOuP94vInJOVxFXAGw15qB42j3EquKRHGSL2bXnrAXvnrhi8RD2FG
MMbXo+07XkplXfc0TQUZ0hczwpv9/8rlIqtpksnIQspZ9ZgYoqHsVd3pAlMAnW5aG+vOT9sciBPI
mzgo/U2+wq1FXmko9+L8IbZ4mkQ7o5HgVHzj3q1l0DcONLB96v4dg8hoDkv4IoTm/Iu0CpQV5Umt
A70zwfgOs9Iik41NU18U8NvcvMuAlTWpHxSITMseKKZ9OohbHW2l9WLN+NWUub0d8yIL7MBlVEeA
+kiWVErNHARaKKITqBqK1PzCCHNgLV2/MeT82AfLukk2Q+o2lRYJbcdEwkurFfrRY2F7AA5fwW2p
7qQpyPPHtbMPW3nv1YLWxElNFwmp/Ho4hrKpm2zN2OsM2eOF1GpHOkPB2DPTrC2sZYhJ2d2m05Pt
mbTrkd/RIsmxjFHt6CGsz0SYvHvJoH0ZAz5YGskEo2X8YGZZ3gi+zeyJwkkRxopKjhlIK3WF5Eca
IDmzrdLBlhGW2f01DoxGgV/PsMHPT8X5WGJnHO57UH1Xd/I99LzbtB8aa1H6UJaPrHT8fh7CIpn3
lfkVe2HGE+6xx3HFVq2b93DQJKIPiqKCC3HFKi3vB2Jj2BdYG4pxvuO6MOPK4lKTv3rsxpcOvjiN
2qC0ZputkjjFqAd2zQ/LHImptL5jTQZ5p9KVeyZXl9at+OPgRH2D6XWnEie11GsaLNUyJXRUh0/2
jI7wlcUqGRYDTN5zmb80jgjMEO573DWwSc90W0Z9109bbs8OKZkKLlEoqQ/8cSQZt6o/zTsV6BCE
VmL6rbM2MW179HUJzX7OVm21TOP0cnziNUwESDF2/FBlpxI5/mA+7+hwrxiFw5nU+BlEstmzJDby
RG6rI2OyiXxXTPEGANWxDRGaPE86wHIiEzfGOpq9BOZOKMZKTS9BfoNccx++xy/j+nJ9qZJ7XiOs
k5QVbtJfX7azsCUpS9dIlifeMokwc2Vav0z5RkQwmOGBzZy7LWz2RNaTrhhRXGp9GjPdLbhOwD2j
z3PHV2NdVP35V+8Ck8/Lx0MCi1TYbttJVazvNSd6ABoPOnvIfTmN/J8d/1TchNZcpx1R7LdY38Do
zmjPbxYnLCY1YgPGpNqi01BCVXnqSrAxfB5TykM0rq2GiDhiLEg3zIc3SrpLOTXCVN/LuCEB8qOh
PnzRgXN1Fd8tcRiUp52kwZJAw2LZt36mQrEpy5DX7+hpFHyEANxIM8W2PEK+q0gM5lemRAhrNcZs
3a5f90v7mlDJ+jwOyiN31gc4w2hhFYeWZVJ9eE1dzD3S69XwN0lnADL30JoujaZsayx+Gnr8o8iC
ha5aI4FY1evZVjdikJ+j9ATUFookal+fBXL9j1g7lmAhmAAwgDMD64ULXxVnbgtaxxq8BVXzCJJH
FqbFP3tIe18/p4b3GgUEMT9r95pIw/A/4TbZehbra+oAjO/JB1QQjHUTraVcq/z+sEmFVln7aHXU
5LuRM3DKK1UaQYUaEst2PTk0JJ3bVJoV7WD6p0z/ySkJPIg5OGQNADjVH/XkyBBHGOh7Wy2n1uJh
NrQUmY5q/L3c9PW71zDmATGuUSbFu6K1GeWXrPH+KEW+HNYLezU1hTibHALt8CpwPSfmCQsutqoh
zresGj5odymE70WZiKDX79L/g1yWt2iyA2BC2qU0c26EYRyQob1NYHBAiOIpkbmDZyZGiaDZivIl
tHl41twl5b9xjkL7r7O5GF/K4IzXQ2p/ie7+zI0vmmWFdZ6En40c1TqUtKEWRjnguULZNTwRigOV
IR+y8S2b9+WmKr2SJBWMKhvpk74YrjErHU4fpTZ4I7q66kLjXgs/rNl3efijwcHZgag1aGVKu1hV
ru45N7V5j/5HoUThErWSL1uC8LIXRpBYtAekMABi4Gb9mNcfEqJv4tEnG6rkovekeSN7JZ58z+1h
HGHLIz7yKAiKRtXqahf+/u8p1/nXI2UJjqT8BvH0LSzyKK405bcSpjdseVcxQnG9DMQwzUKoI/go
iUciA5MjSYm7KKptiF9249CqKa0Yef7GViffQPpMibVVnVk1WIbUholJhVGO7A1TuybPnpLA82lq
AQFStLr/7x2RYTBUQkDq1mtmzVT/1lfIVwz6e0gRmcBUuRjvMc/Y05AyrCFiv6yCmhZas9jg3hAN
KOBlhFIv9sYyPRl3WL4pXfRwS5HNpf/+Z05GFCdMdRBxDFx+S7vocFBXsQgJE1vjxiuIAr1Kq1xd
UXTgKRYMdTfO/xJxKplaLjwD/slkqDC+2a1WHdeaFQktwDU3teOwI1v3+xLQHn3FiVL8XQz31zNh
HxfLVUksknY1COIgvjh3hFf+vxykG6+hZZL6O7Pu/v/xuVQKuVOuJfqflJUUaGZQVH/4MXsb3EN6
IUU68dNLBex1/PRiH7f1iqtzasgoiS8fC87AG301Q0opUHz0jYwHUG64e0emkI2FkuxnxVewz6wJ
bbXufiF4rh0zm3FGnevF5T9KNvYdwfOe/C7K3sPHQezqYk6/42LJ3A3mQC5PgiedZNExxYCSxzqf
25XAHKtlVJQX8Z+c+CIbu8xcDWH+969Se/mwb7xYyXcCokgJ/uGHL2DBh+5+YNfWVFGw3FNC+2IU
ylw/+08u0yV752faCZDqIRdniQLV7SUv3jXzia3ObCFlF5fLNgFwWlDzcnmDHt6Uv6y4aT3Y8ASr
LLh1zPvqHm1PJmPFjcCXlVcgMtepl9uStpD/Kk2kqF9ZMpJCfR16a3MhhjgDDv3wiFKGfIg02I4r
e45X1JVXswUQ0aV+yy6jXbIhF9eojTEzzRkt7l47Dnx+jGbQIICNBN5/PiDqkKg3hI+L8L+J64x9
aO5cBaeRJbDsT3tJwdOp1jx/zeiVwQwQoCne4N7i1leLJ0WU/DXXf/J+vAPlMHQAlnztX1z4Wka8
larKa4+DuH67kO5BeFBN6O/jDcd2i1H7OhqWH5L/MkI9XvFUFWlcyqgeD1ed2S889xvkT9Prcxp5
THF3C0YyRhKK2rNgLU7sY3eBb2/jHqRLN91HnUUirm9omjHDfoaHzCRs/bilweaFoLjZuDWqexXw
VS0PXn0FK9GjQ47vStN48DNkLP5tHBWkeXk0239eSGv5TNXUTAl38NGvcoOh3GKqFelmbrd0R9HA
MObPncgWnlTtQV2OaiN8RSmXHtd77sLrDfYTI6HHtxtPSH2xSBj3NByO47riNY/V5UmppoQQcljA
inewWCSxUk7nAucLcmeUWUzjMcib1fnAMynjPhTSr+CGX191alVOH8D8BiSRIlVE1rGKcuMpOrbN
VCi46KI9wbk9AnepO+q+wUOSDX9tbWbnsDfrqjTukcO7HGSXLw+8jfPlfAEjwxyiLVGdFHbsK6kL
NuTPAI1uD6jiS3jl1ojuEnjbZsEyjtc+DIa7r8HzAj3ToGet3ohstkEGNmwr//eFiK78EMPMiZ+y
Ep/GQ41/w+yG4ypPIi/EylMij9K/KG4EfkMCCHIFp2VmeOhBQKGNo2CgrP89Ph1LRsbRGT9or/xJ
xWnbiDkJV4fvzRMFa63Z1JQFc4m2LlSchBN4YX8lNr+Zb9fe6OJCnUmHEpLDP24wA0vSPJPqm+Qp
RZ2wfQEnGsa9wvUSRWV/vPT5e8waR7Lf/6qtePpds/SydNMKsg79rMwPAM8L3np6ranx9aYKhAo+
MSvKSqXmj0lsrfgjViMQ7SgSSkyE5HM4Qz5bd22tQDeAYxOBLkIJeuLiBarHmDyhclwfQTgDKDSO
8T6VASSsxA5mc1MvxIDaIqiU+Zqlbnk6eCJt7qCrv0KIlUeqOBZLv/kLuajerRUJt8VU1vPPL5kA
WKWXOP0okbz8DCPDmf18aEAHGB8N//u+OAdpSKk9bn0sbENsETFaD7UoKezd9JGtIRS0Sp4O3F0i
+uSJIBESEv+FtAs7+aGfnnqwIYiOaVhbHpTilawnYJ4V0xaDD9NkoBEYE0BsBK+Yti3/zTk7J8+9
2/tBpYIBjh3uJEQkNVXwHalxehZdgFYvzw+e82aOSILHDlJEhF78Ahmonzc9tbkhmFcFnyzfbcqp
Bl4jpNCdJ+g8bJPCJfGCheAcN44wnHrw9I1mJcsMYdoU7Rcrd6PytcctptqaflDDUv2BxhqczFv1
/FmhrZGOJbVtscvVBp3ylNw91RRHDrHb8mYVvFnzUUXvrzQQ2gIEI9a06Fy8CHZ0GGJvjYcM1zd4
/7T4GqnQBQacQzyTcPlr45YxXEzeegpJp/UbptymYBki9nfmefMjKv/G1yJadLTYXKvJdPINpXcg
YM6Z06JMgu99f/wSuwEKh53WuHGbPvUsC7fUEBWENJxoQ5cmHx/KfLqfGNDPBzk48KssWiqTg+Vd
ilN8rCDD0SuRe697VJ6clb2BT81uqTEOrv7RTDLhytFYRdRA6ddDBdvjHlPsdmBSU+6iR+8IbToM
Zf8f2jrX5obK9nkeW4ahAJ7uRJ8elhZdY+c/gop7okHZ6F6xocuI3UBmPU/U/UZvR7phFS04JCM3
zACZoOa07adgamM3K8YWyh3GWoW4cU9UE3oXhAfa95VvmR+R1aH1p2HhnwZIjwndNzg6NOYEl4GR
isyR0ykX+vmdrmWUiwxrK9q3UhUM0vwbbdEdKsx6fQgEX271qMq9NWIYy4orraTWsDt52nxjSUjA
VxMlZogByOLjVyXS1YoPK4mdlRu7zfvSFWvVRy35/cXDaAJhqWZ/7sZkqC0Qi7/7tN4RQyduB1ag
CPzYw1RXSXXpIz1MKd1VWLeU1i39lJ/+VF+I0FSI/TTzdxdPjkFT5uUmr5PndSfDRUff6Gh1DNQN
4/dBO0mRxRpodVs5gFhpuMu1W8ni6pO3Llri/cLuDErCYldH4jTu6OAoYFXn5Lxaznp7NHAuVBE2
1ewfWnsHP/Gq89Tkm961U2z8k9WwrQlU+gyv+fyD9xLyVtshrqkw/H+nssM9TWE4Mn32OfTxufik
kBqLlpC73qoJ0i6M7NpjTp0xoPVmgYEXUe/jzuSEXUsxwCMFHSjsplXGWJNlV6v99/TBdhkSwPpl
Fzqk0g6kglFr/QiqKmiVvVkbeqkWzXylHXzpM4ACD86J0FTzoox7RxEzF69e0Nr6hznqkfXs0FmB
HG29Rk6sFEydcoVfmEj0hRYjdVlYCEu65xiXBMx9k91wNDPJkPvAJDftg4jr965cah/CwF878fmx
7JQfjrgVZQtaaicPiaiBZSQEmmf85gghpof+grWff+eZQ1l/dMfPziP26inDPEupnnfqylJMP9BG
H4IZTXAVWRjtuwfBVEM+MD4krRQE5yYy24AFeBby1LsJ1ra5cmRL2797Odlwj89Pr33R32zzCcj4
dN8OBsEMfp+8bx5WbC4w9QB7yIie91kVOGOhRgm/UTtLv7Ij/wW8wMLxUzN4sm+NSPIfUNWxrxx9
URWcC5uaVT5OA4yAiXqECimqPF2iQTDoGXcxeyp3cNYaseOHGFMS5r4d0GhquCzcShx9SLHQ5JsT
HGSPbJI7PrAPicXQsmhKCJO/p0DShk3F7Obq1MauKngvRh4bjw8oYnPLKgloZ98aQF3LnE0bP4ph
phcAPRbW3ykUOPImVQtkLpBf9g/oqiN6IVhVes9QHggJ+pc1hzxdSnqXKf7XfUb/xyDMWdi7hEkP
PlqMXwHZtbAdBalWmBzkR2+01XLLESg5j9xSYTn3BAt/2LT7rOcXNYgEUaFNlBxkFi7SXLDRQO9g
wa+Cof2X9OevCyIqkaUrz8n9nSGUUJRk8r09iCWzoOlrHlowxBBv5uZKRHg79tavuf6IWRb5pJoi
VlZK2St4JV3TlG7On4X5ZOdVbgO8FGeF6oJ/ZXeptFeylh2LJaL435HbDXA4L0el7OBPAsjrwMZG
BxXDIX96Cms9g9u4QxLUy/s686Lh3eJ97Os4SZIKtdZPrQRXu/zQeb4ytLtlrrj7kQGdL3eFqGdk
NHGO95BUbkrTHeVJQeHmr6YZD8R799kWhRzRd2l7epzwJB9yjVhQNZIGh/WUIgaJu+vrY9eBLKX5
Px+2dnTvdg/+f7HSLbGe5cUIvgFeT5u4KLxF3pFHoDYw+EA5JbooaATaX7uwNSg5gYF4IiT3mn13
PMyJEl66aZ3UN/4slP7f4j3PL5DxpQF2VtjKdrp/a7CNjuh+SLOs1RYZLWy7wzUbwH43N31/8Wez
q+o5PFLcrAcY1x2WrJxsnNsuoHUlOT60+hFzDdEuEkYAl52PkRS2uaCLqTtiOHTCRoaquS71JCHH
DqfebMCscT7CXFK95q/vOSHe3Z0PaQ3VOUPoA1wiRtKinHZJ79Kc0c8XWXPcbdKxlYBCloQ8eoxZ
ELmZ9Hr1B5U4eAeFCOJfO1YHXu2iK5nT3ZOB3f9yC9+MMd1z7jcmi0W9woZRBK296j4U/CnFDUqu
k6dmz1C8p6G3oUhOqQ18iCcziS899pgqFLSQcQbbPcEA5tPkYkVBBnTnwGGLHKP91D0yVytoC3U0
3AD38k8py8JnZi97Hs0zPgYafSTD2c42K4Lu6hblIDM696aBDycNF36hmdl/v0TiGFlQXQCKH1MY
YbY0QEglvU9TP2I6a8WSzR8xGlqacICBkUrmwHBfuiv4Nr2csScYLdx/uBYDYCLB2j85FrlRbWTI
eKXZyaB5NH2+hebhcObgO5RD1ozIxU3YtwNxivspQSurrx1SXqRW4MN2vvb8U9+MS0PsbLIuTXDK
GYRnesKRUfwrv1oCmNnGc8DXuSv5kbAYdeUP2tByMcSm8opzPqtG8JlsGQewipOrpSMKrb2LcC2E
glEZHvZ44q++yQEoGQ7jlMgcoQx7Jf7MUNRhwkauPcissdeLgynxdrUdWl8oxP6UU2v+K4qUmRCL
7fYV18aZ+arVpg3HL9KR5HZC9hgID+1ZupPaL6XBU7SboRt+nqp/BtxeAy9fXGMvF+r1M0g15VBA
yckyAEUfNBiK3GH9mVzpE8W57VpqwORyzss/pbIr4lbMBC+IJfKAPcw2xodDzC8gqA3BbMpK9L6Q
grNcARzVIwRwSGvxgcFNQLqXSq24e/2umf1/is91RgziVQ2zkt2E1Dp0AYwn5wq9eL0LU0xXsrRW
kiK8ifbidtBAuEK9B1XJsCvCzrcIlJouU+nGxPWqV/sGBRujVosyjPa9tma+PGEnVbIlHRh/OGS/
Dbi9iF4jbV/14ARll1JM0UU4yXSa00MocHaAu3mNPsfSV/KklSnaF9fS3qmMLMIDbofN1a3vA6l3
xh7XZy9RjAS5RFkAzciu7VDOum3xNAyyw+fl5+5QDKbqt7fp01I6JcedckvCTE55aCeQTEYRFpeh
XRGxO2NJoWrvA/ku1dHEj06RDbBwmyFyhqVfOyAhgKmli7a1cfBW/SZqEZPgC1V01ujharlxQGs3
LfW3eYnsQA+pw2SlrgnMhTjixgGspm41hKGIKaeosjuLNfrvNG6fFk1hkwQBTneq7dncFXWHweKF
l/ynWZUOdWS8zj/+HrYHEUQs087BZb2AwYcw5Lr/XyeW+CaYTYrX7/Jq8nH0QbWlx6WyELbrrpV/
1MHxxdgbVkucCfT8Lh/p+YZ4VZAaaqfSyGRbIrivkrLmHBZCYl5OPD/CsbvEwqFQMwsp4E1KYhvf
G8ZMqusCnwOT+h2dN9n0kA2D+U2tkjfSqqKdV44Xrxr90BhKqVcr2elY0ows8BjILdEwbkT74Orn
VUVM6Ll/SngOZMb4sbmtrN6wimLwuXt/8c+GhpGlFtlhQi0DFalzkVCve4H4W4rDModoNf2uYZYK
uVOfEVM8N8gjuxSu5VdXHSwkx1H0arOjQxuFNeCxLeVVpxKMeBYjOvaLNjHDz0V/PDqH4S5zZkM+
yXQOksOGlZVzTJQIjmEuhYYLgVHwDaBEurcBnFWUdam3H7EbO3ZEQ9pCzu+ZOjW0k13zporGp9aR
jLE0YzGQFpVrwBugZdpIlWdwmO1jX5jsjysTrpi/4zZFTomiVkb+GYqNwhs0Fh99AcHhIanBm+0M
I1o87cO2Jes3cUcH+79Ew5PcnDFL7oAa35XmaNAofh0+wpzt6OAPfKfXDH6k9A9pAO5VZJYVvWJe
hvTlUrF5y66e6BcPzWgX5y8rhq8hQpCnd6WKY1gf2JhvbMroxY+LIazUQS4WZkeJPPB2U9qZrXML
kC1C8PauU+icv3jfszcx3NEyhNDPJw6ml0o8w5CnmGrHNr2fpTVN4n2i2PjBvmjS7ffnw69vJdnf
rd2uqZsq9NJEg0u/Fcx0xeB+jjqky52HLvklzINdwSL+2WLMr6H6YkrM2YOMux6QWOlde2WBg65Q
7gl+UcDR9kUV/VH499vWNLK2Msiop3VWgIkSB80BSFkjUMbXs7mlrdSYAFe05t/hdxRipO7ovTxb
76LE498xfC9h5iolFDzKVjjZWXBqBiSUK+Zifnpk10izyZ1hsCyL9ST/hVFv5YYCWexx9MCapiMB
EougOCR09+D08r1vaA10yDh6LUymaYQgNjoNGdHLDqd7U+9Jk+YqBxa3L8XBFlaV1N0DYULRv9GN
cs2SwOqsP07/V+0cP4/il2ldvB4jQvWIaLliVHQp+zfAd5csC9c1gp57Pgo6dTbYmWgN6pppXXVy
7ODuSMXOMM4HOrJwm/aHRtR2xiJXMn/XqVz3BfcC8J9RNYyyJkUgKdW/no7PMljUBShh3a4If09m
o1dr/K75A3fPF49idkGIqTe27MB3RRERlTlo+FMZNV06kNN9mX02TrWNSo5jdSAnu8UnV5faYDTL
Yrpro4iQ2bpmB5HTHLCCqIuXm4iPiMPfUbiF89GE+3ePZNmHZxjODe+LVgDo/Ge7/jACVvfXhlSK
mjKOziUUEeLXxXVXRUIEqmlDZgWfEG0bLLGF367TC0M8Rb2WQDw7AOzjnnvFJQcYYn6NEBc+dSsB
0zv8xC99TBSUXun9JR4oBL/91KLdfe8vkz2qRtVR11nfUyMMg+lwE19KaFO5NpAuIcZUDO2/Wnkj
TNIO8qQp/+45HUvBX7hs+JJ5bkL+zd2D1YDnzD9HShTfo4nB313o9jF3Q0lrUM3C/5zHbGnpRjQ1
gZx0MWhJTXsCkMM0gX+/5Y5+NiBzrRki5wvMOBwWNhtAi77SD4CENmNdDXNBRqqkBdkLUGOseybi
/BUo8eH49hCMX9TM0auooLOwLIV+1YJjxhxoKB5nuUSOfPYeaWl827PwhE19hpM/aiSPHEhFPFES
tv8fbLMoCi6InOyO0Rr+nvz1gw10Ekp82RiR++yZ6PRwFSfSjO9B4wp3OL+KmzbMrJpC0DC1aN3I
F0sm3U5/a+FRWRCd2MGpwIR6U+xCn/qTqsDrFRobGL3sbuY3EQrXUp+THvki9c6jtig02i6RnLUj
GvNvq5bT669mm/HPU+JAFDlNQP8ERRWFwPmN+1ojbrbsD/FFMut72vd47ezq795Dlw1epgDP/Etk
YGTPuvRSMYpUbOjvBqRnHaMIrcvH2FP80ngSdppR1NO2QdzgGotaZ8WO49p0pBVee534fc7M0o1O
yZ5owqfEFBSgPNoDAqCEgjhqg+iMDPfinVeH08hqWapO71J7EVPgc8cNgPXxMkdXrtCh02Y516Vk
aVDuq3L/H8V1MqVVZh5ie9prgnl6ICeG+zamoCSCJOoLa+jcP04a16HaRMGrIycbCgccOHThkg/g
LCehBYxyDRBu5AxqL1DUxAzzvzuXNTZIKywXa8GHnQEmCejqIF/dNXite66937JGaqd4Amii6kV7
Nck06pDFXxIlGgnEZ5WR3Ee4P0x73JZ0neMqplsna79J4MeyHgSamsptIOK84KQkbU4fgYkHlfHX
j0eHtVNqrGfXFd9/nJmpKzRCuAGikIdXnYHkz6BcivvDDhZ08eORxKnApYxEeoZTXrd4nS+lXmfE
tLIYPSY/tQlSe1Ap4Pj4USD4BbXNGp7dikxk/YK00NAWLA2YpefL4MqHnqkd/oPNEKS/ZOwkd69r
Vn/r5hJ05jVkRQWylA3dYLFmCnH8QetiZaThApaEjhXwQhf/w+IpJl7pYcel3/WkNZpyKJ3Kkig1
LiuaHziO71bPj6RRVmD0JLOxT1PCzM/PtZO1X7IsOO8HKLzPUhNOnFl8Kjkt9/ZcOc3yLJsqJjhE
XmFmI0qeigzx+yMgqylU0hyo7M3uROosTSzfx0Xc2AHsz11gIJo1RmIBghk2RDA3gHqdyAFgwsr/
bzgKejhWmJcG0aeRmJQ08j1fzYwT6R0oluzppXryxbsaITlvY6m56qSz5XBo1iQhuYXPrcAYQjDC
y8Iyx/Y/SqA1RmFQ8JwwMIt5Du5nTk2J32QEA58Wai1qprZkNmiAHkxbNyWyGncs6HQVqnsFHmO2
/vTdZmQJUbQ6DaRcGxt/WYtJHd0RxOlD8qln4vGFyh8Xz0g10RhgnvCD2L93ERS+ynaUmwd2oLxN
+EaFqYh8Y/6TD3Jj6VmmLzyHtMrgSwZvvwBVIOY8wU3Qoo2jpeptnC+0bit/a2tjLCGYR6drwWol
O6RppY9qK7AVZbtnnhQI368qFVYSaIaqtLUG8I4+C4zgidz1mz9eqiFI94Fwon1HoHdK/k7Rg9Xu
u7+bioQnCNRQ6ochzje8PLPm/fcnnL4ZFqkX5W1taK/1Yduq8bMDRnMgejrpNGfhwgYJQPAi3YVG
9t1G32wAPxO6bj8PZjgDImMpK83vE/xWLdatNPvlAWQkhfnRJ4x9C5GwB7lcDU0YPqSVRAuUeaR8
jykVihrpjWCJiSB2cPmCOhoeglU76djEssHyEC3CeV7v8vbjb0RRO3PQXUCwqGFtLMrC2OzB33oR
e7EWnry43AvgAx6x+SDZWc1L12TVg872WE+8BJo3brZfCeEvocfcLmh32s1Y5mXF5Psb8/1PeNUY
AGnr4jFafImzHLqnUBs28GB8YLlm5DCACcUCjGfhXiTBj/beG9YEFRrar5aCSbRCxEIKpw0cZj1n
3qycALIXbnESNOrRLcABrSmcUwADZtpZtDjzsU7gLNgippQRF+J/sJSWktfqcNHvYOAcBNoyvRnX
msJV6uj3pIpOPVoj660TOvdiHDiksdDlyfg2HgUJP+uaPURIG8SZ1ljOMQAU21aXdqNUdLunNm88
t7tw1JiGtivaInD4+AG6iR3emD/i+ev9GFc5bPSvOOT/ODCW1UTgUUBVlxkXkF0Ze0a7JBBXzcwr
coZMIzSMgChIsGfO8Ga9OtdlE4L7raOMoANwRIT106so5j3ASnogr6CA6hUenLyGI1RCRMYUWTq6
1xyYZf/asXwZoqARLObW755GDkQK5x9dvM7Nwio6YPfx/1QHv6l8eq8BolYb21WvmOHFijOXiMGB
F97GyfxSdfmpvc04T1NqooPcyHHyRrel01mhg51tjqMxehWzFPCZ0eeig00QvExGVHBpUUCywskX
SMztV47QR/lmnv1NnBiHLFFQveVy/HMEjRbC2IzpEf1O34+TmDnQpsuz6j/za55O7jS9oncxzTSb
hVUbKQF3UTB2pgWQIabd/AXxGoMHDYYFTr6LbYDYAGYNHqYjuePiCx1lyp9+VdtfnBKUpqXyK4Hf
i7465NGGk4OpACT6CJMV+0Rd/RJFbxEOWyfSzHFB/N2mAF0eNLuUesrUaJwH0p584KB+wlP2pQNx
Xx43KLW0ANu24oHHCfkHM1EOF3N+BGlcQviU1gk5/oQN86viGUEdk9IBAvLA4ky4RQ8KuKp9wxkM
XoISf7pB2EyUkAxqUISOG+WEMMJyI3aZeRBxDuLkqd7HL3rpzc3yfEH0sm9sGbx3OvDXaPDAmO0F
Jv3SPapN0tgv+NZJUFIRneiYIUTOcGkTHShBy8L3+OJ2ts9M7ivodPTto37NOOYgdUM6xK4urQ1F
zcnu8H+oThaC0YiV8pFwZYIDWxAXNSNtWou1sF6/9AmDhcSQKVcr40SdniEpeTbBTcaqYTbEZ3Ox
C8JnjxQxNxJiaFC8JyPzb2wM728+kTeyne3Mjr2pa6eM58Pd1yZtARJbZWGr4mVd2LdQxwNzN90O
nnB3gPM+wd1ln/dcP+9om/RcwsOBNk1LhOjfoKoWRi909Ax2z8f+pkIiW4+4TlZ9QjZ8cuPaJCiE
aWaENXjiMziGt6e83aM/qfGlxOGVbwlUY8kx7uQ/hBG+WayQDk28+jFxV0nh4ByEe6I35emXPYWf
WlMdo+XOAfOllmj4pU9BACJcikaZtV+LBWQ6vhiMF8sBCruxdkWfF8uANx9FZbq837bpBQlBkwDK
8l8ulhO6GMwa8QsRMeBwz696UNkzZF6mC+kilG6XdoxURv47Jk/joOpoG//O+cNxutUQEY7swZuV
QqKpsROaoraceAkKzXE9yCVqtbmFB1ukMeRrZutr94SK3SF9uYSWNUg1uU+kHG1bog5XiotsG9eX
cSnLWdQeE3Htsxx+tUy5CTt560Dl/ec2z4A60I2K+IbtwToYhdEpdi+cjYjqJ4kAisi2D6NDlBSS
JKW8/Gtol0cOUStoV6mnQzCJ+RU/L9JjeGBlL6LiJq6/53fpPQOhsoIARPXzrSdCRRGvZo7g1lPd
lMXnGHqRnxaQQVOaLK+FN1D6JJU4+nAoApbMl3kvDhobmcsgyCrfceedWL/RSRh2woqtH8krTs9t
pl9xI2qRMqQ0GXqwy2wI2izQQyJKh11FMpWjekYXd/xJBssGYGamMwpU3yr3CexIhvTKB3BL/yfi
CrcDPCYTP4/5A47kHDVilVh+YZT2gA5K40KKD3OGpZKdkWQe3X8xluwkIQ424kY+7Baa445GlDqS
egkBBVy2y4aVReHQeu3x7/pfDlvysnCMgbkMpyvNAQP87iQpk6VuqSg+beS3Xia5aarfeWTFXR5N
piKEf4xb6aV+I+ZznF16QrajvIUqEK2E0cjAAHqgOyHz1N6SeGObthsOK3Xn+UG+fiaT2og+8W/9
wD+kBASeYklqknwPcz/RxEwVRIrWvul1KnBA+P4Ur+/iyKNSR0pwoqinofa2kKtQiP21LK3V/X4F
EMo9sO1MW9YyEh27RmZfgLURFOEQByk5FPdniWLtIUZkchLSEkQ4VtTptA1K9yNknQ6V5TrunPdP
Gby3Lgup+pU2AmvDAEO+P3pA548ooTj1e11SdqIKSH4mbDV0Xk6oyCO0tD0j6ZuxZmnnJpM6lFHP
HAKBs857Sb9rw5xmrRHnA3bNDIE3Ls7vvc2XbpPNWK5aqP8ARIrQ6AXEefMbItuUMtqIutaN18ot
HNHqT6dJDbusv1h+rEf721JNKTbpLZzRbqDvIAhTmPLsPOkgWUeC43Ti5qgavjUERQbAi0AtUYRu
thdZOQeN4TSg+Nth81mLfgxREax3EpezxaipTE9PfR0iILZZLp2nr1GKws9iojbL0c1yAix1GQmT
DqSc1qDoXT8oEcIfg1X21dzpMHxJVhHOeBLPMV50Discl2FI/fqQc9IVQyZfKkebQWS2wmyVK2ER
T1fv1sxzDXdF2CxlMwkqJIJ0eLOJBLngKgHJpLw6G2Jt5+rQUgfBjeJwsF4wwuGzUOSBCMxB52Bs
SOD4wdZIGE1YDP917gTTOthZcB4N+uF++3I7YXFHVU6HH5b3hLVF7KQme8Do/Za3UEPi+S8yB92K
ltgnzvFXvvN2zJegLI7E2nYEpAkCQottCAX+X6GT4jpBFWg8+YvgngU9NKjIruWMPTxPsLEpVzQS
AC2fE6gpxzzwAH34rTthDzbMLbLRJlov93pxfItWyZJQmgfGPAXtzIIyGuFNDcZYPswL+BmptF7U
hKSETum0HgybIBOUO4DyPQhAqczvcE0Xg0KLkRf34NuWauBUs+b6V5yxBceDhmtURQIszZlFPN8o
1ogqFz4bhcccdxHJjM0fplMAk/dy0+sULYlhcVO+savsz098l3l8U0CcUfM1JRIuRcGG4SS/TGUy
grQhz+/sknOeb6WWGta62NJTo3bWSDwW/IdDIixJnZMoEmWZsYTB5M555ZPfemtir8ibECQ/F5w0
b9HfAJt/LyASxjYXYjj4CLevZkV/EQsYrA/xoBJl01xseFEIpfNqkclresXUHzCPXovb2nVvymWf
uHRcDGBoqM9Nvzwop9DoHaqMnbagPjGfn3VdcPQ6QeeR/R1/7xPNjW8yZmptSmlG9JCt6bR074G/
5nIDjpVBYI4BbLZkCkBilqORqFhugNq62JTASuQDxIu5tFGjD5aLes4WgMLYtg7F8R80P2ekQ1GY
wb+DpbvmZDbpdAFTvtWQSZFfas8mzjEP5EdXmGq9M2Kt3YlsELCOTzRTQjIFav1aumnFWvYkTIMx
tf1ZsdM7ERG3SUTkoRIXXJCxqjDiMYXwcWI5Iqr3MKUYy28HXryu8pXI9vbnhdK+zJbdpYnfS5GY
wTwp3JpmN5d99gGkvYLNqW7VhOrmznRXFSJd9hbQmuojWLyxW3HLX9FRktM3p3Q+n5ktOhj9BQ1P
tryCFedjr4mcVAaqL9DsFalHcKaK4awcbKy1CL6tq/mfb3ozP/9ZCiysb67WLLEBEPURoPU4LfdW
crU5/8ImI6cJfON5Uw1y/+ngl0aSXDIaoK87zhTg73pzGpSvvSWCxSq6ag1Dz1uVW+UnPbW5ot0k
LfJlf8Qad8asgi9L7i5xDq6s8oWx7Yx51MC87+66VsLQG6EYxjlpu8I9/oOjRQWY3zmC5nuUgwhE
Xy5ww1CoBIS1fwJt1TE9k+Z1p9ju4Vp+ShbD84ooJVJinYEW/3yH9KOTlvSlIfrOTQC8EMgWBj+U
OKXD2YEqfOfvimjIErYV/2GJ1QmfpAALEr9k19OYcg2mh9yY4P7OfRTkBeoTZCHEccCVnsqtFWkt
3Jqrk39H36PdjXwWeHE9R/rT2LaHDTwQx32/UbiQbrb3WFPS+AP56xZVDPuB819Q8MRtvP6+8HT+
dgpKRxKCWPGiba43dwyyxJ7IrtezgIREy9RUjSQ8hMmMqzYjBbFpAbm+trPHDLkmwOBFFcTYGHzn
blpQ9wzGXB8vlBXLocYR0jt1k/c1OQh/lGaxw82FUFc9hJD45ONhsw2NtMu+Z8kTT17vC3D3n0Sv
e6cNaJrKLTZw+gIJL+oem+K7osNzm923KVbrPUz3PoLB2nvJW0pA/6PhRXpNFTE2YFyDF9IpSohb
LHFpS9sBHIvj4spqcTTsZJMhi40Ti6dGws+ZK1gloPyo9ZKcFbDxB346eXZpvPTSY9Jf7DPg8GXR
AnVZEUu72qYwSgsNOmwaaYbo6TQKrGJTAvGvnBx/2xfM/qNWysdnypkERqu15H+KLw58/uiZvViC
gUmsU4heiXwgzNy8Qjjhi4Ywh+sRxI2ZtLN34uJ6XMEEPYePqUj5v7iu48NRV5g7mXufgxIcIJCk
cQQJ241ZLzBQRJyf4IUHPutMX8TzfOyjV5qcLwd2pf8gkK32MFiw1ZfolRvx7jc8QW0EACTRZR3U
jriyWMo+s9JRIrUR65FUSgbgCGWW8aA47Td1HRyYvH8OHYSCZZFn2Z5xgOEYDkmwWAFFWV8vI4xS
3Pkzp9URkpc+JpNQuEHzQ1v/L+y+tctlAK0WQMV6x6j+eTxFS9bY0h+JnVrKZtqvdYKljZ9tHz72
kx1aMivtJcWYqUcHaZ2Vioa1VdFLkBkeSbebNemdas+qo450zWk044LJKoxlF0C92q4N+ahVTHnT
9TjsKnM8LylEBIdYvfmcl09m2MScKYKsqeCb4I/l4e5JeOkdgi4hQkufrtOXZ4YG7wpVDSxg99KN
nGKEICX6Xa9c2Y814c4/BVRFyDtrwdckFgbPqaQyXaRl4pGNJqPpe9Qp2gi/h4yuqwrVqEp7aHsZ
L4RI37Uz8KbAqwazN91TLi0AK7Nvim3ZvcehSeLJ7Geg8BCSK2H8hZeRXyxKQG+N13R0rkbsgvVh
ejmimH4Xp5asZxVpbrNKNVVFWiL4QBHHZM4PebMQySC50jIqHr8N5jkPBf79s3/W+mwejuH+ZRtE
JfYHvQW2zenOMOwDpDZcWoAwVBALYUYoLuF/aupVYaJDMNNPOCdWmgLkxGluPc5u6/8NuVy+c5Y2
cmOd1stMFy2nGw28aqZMFBdRLym1VQ8qQ90joR8M+nVWENG9S0QF1PEM+ics7033W0xqLKMm6EM1
2m/BpvWFivn3kv3yML6euOrIpWF6n8FSjOJSui5uwKP88yK3nY2moxXV6fipYFR6FMHZpVKucIA3
nDGCv4bNFn5RkytxKepdsH61aCt2cGfl0tAw5q1l1qZoHN87mHNKYW8Di7AjN7GsNluP884z/uwY
blBa1q8PigHGDilX+11LXCRFca7AqH/KQ43LruvmyDlDtDZn+x3308TtYXrygvjYbqPL1kjMi6kU
Tmw8clsdULiyqdaRflX48+emTPDwoaz/7rx53nODdLLi81I5fDuythp6JYHfgl2I03q/0mk6uynC
XkpV65pzUDHdy2y8Bwe7uAc18vyWXCIQuq1C/TdlBUI3p8fJuCL8ICoPc5lvhPFqWdnk7mkqALlD
iv0YAiPWn9tNKuEI39TSMmMacCXhtRD1J0Z592zaXey30x+FIaqgahc/yAmd1ZckKZJR2zKyO/tI
2CYAYFrEUzgfW1V+S3htnmz21WRo5w1cwCCUKoHWIOJkq5q8fQYrAplGMpDH6n5ipnmzq3A9NLn8
QKfFIHzM804JBKiR4mBuupdPgy6d54AcrM2O/gEg/R2aii9X3xoHglt/+DD0z3ED18fhnQhFQ1eH
s2Bswl3Kl2FxmibDyzY0Lxuo3kkqUzRtBK3vcB1pIaRGe7bG/0F95Ec4uf2j9OTFM0IrP4PO1HS0
igpDf/TG5olkgEObGTSwqtSbED2oCPaEnx/eNWIB2h5/58rH+s98xTX+uSAi1lNNgrQLFOGfGdmC
Nd6bPKFwaYYwZ7nVTw8I8nnjzx0gw6Hqb+N0opZhYC1ryS0qWN3alUAUK94CBK7ButTYlkPudVNg
LN53P0r2Qhbs2WIJMcb9tA0EBv4SyAKDys483S3IzZ1MixPRWyFpyz/GYaYCngTAAZeXmYl2+uSh
MvQWUlcARbxsEgREHTzfssR8hi0TSMFeaUydhMJJfGCrXVEIXKKYvZm4uHoeK1DsWwl/W0DlgsjH
6QewRbj+3jnlkFD6NSC2vCu7ElbtgBsxyuH4vn7168DLl1T4VQ2Hzpk4MLxztfpB7bN8CoRDzn+m
H9mtMv6SfT0sKaDOHsupAZMKxTTq9Ipa4TLj7XACSPLjB2jle7EPG9tB/IE2Kupn+iX3UyfJKcGB
XgXu9dCNerhf+C9464TBonV8oZJNMgTSEwxQmyxU9Bd8pgoQJ3hYD89TPXKUDahkwxmHEAMGBEqx
9rFgx8QEm70PvWyQdP+OeZVAOX4BqY+EK6wE57KeMNGLqiIFq+2yEL+B08jnxbVq832Pm/veB0Oj
Y2duJuyrlHzYEVqFwmPqRuNcZyaCxBmz1wa7WlFYX2k3xlxElrLWSAmf0uzTbax9IwWZqUC4rPc7
bBT4LLurtX/J6x2iMN53a6bvJV5jCWHtC9/OKTi+eIdhq6bpJ7ENI0ylWXB1L8eeyd5n+wOb/b7u
rllgAB49r8N2Cujnb3ztbiSKjWPCBervBjjVnhy4uxpZe2DhZmLnS7Lp0tMw3O8IN7oFPK7zNd0G
PDGimVJxblA39VzYplt/m8nR2AasiVYLS08QC4eVj9NDTA2Cqak5yUII1gdmHeqAoKiF4MhvRI0r
HBpy90X47OAEpVy22dJKfPRsH3DhGNqpyP2xJQ0cGpaMfzM0952hqbtjp/rzqYlzWxUDJLRLLXEq
K62NYhIbwoQ+GG49IUkHvWt3Bh1h5sEX6IjiwX44EpP54usn9kMDX4sg4mkPnu1G5tQEMeCp8uHo
AoFPaj6w/DesXc0NgXz6vofDdDhayYETZMbzTBEtKS7cY7jgGTIPM8tLy4oNzuKDUUsFYhdUIH7j
yQZL6FTnk0Z/oLLIt/NBlbdgA5EdBLiWJpcHhkb6nJiuEEmJLiY1wHm2CsjjKnILsIyosq4fV0AJ
qj3gmJWgyIrLjHc9OLVLtcvB/MT/AB+H4apelc08WCxE0tqEiC0Iwb+dO2ISndW90TnxkqX53szq
a9b6ddQtCXCLsBOrV24CopI3RN4dF3uDmyMq0ZDB/korSylKF7vJqLU2GnsLlyJ8oYvHdXaXTYmC
Fq1uwEa7HxfGs6Koi4hR5rD4kXj5nxIl4o6m4wg4ICovEz5gHf21PKwDP27pSF3c17J6ItL3PvFi
LQGN2XAMI1b7iz6Hs7iFv/6My3H87HTM0NzoC3lEAIqFiNgYdiPr3qvcnieo3AZzw/ccv5r1HqPP
KwzOSkeST9rVmS7Ogp/jWXMheUZT4rgXABga5OkGkUPgc0iPjEm3RaSoG/AWlf9JhHNZC4EoaC1I
keGSzd/0f/C1JqhGkaA2UDnzYrDiKo79bC327lz/fwHNHaGBzsiDoDVQzoOq2n7Bto9cdUe+dpof
c1BggiYgXVsbYgNBEroZp/gwFor9CcFKDLT9UmP0oA2GDNr+fHrGibjNbk532ufRM51tMCuNnJXx
du1sb9Cg0nAYvsKhT8IOlbAYZ5gijLamuOF5w1C+BqFfHP8m3lMRvAj9BfCANYlN7rdJmr+NcGac
SP0LBSSuv/uUaYMW77TL3pkodV9v/kboBDL7CBYgxsvU18HUdoQT6ohfOA7dMMvePMfwGBUENF0Z
lBBtRrslsSr4mJ0cLROImvQROEkup8bWyJ8syDEjt/gVMpcnyIK18V+sSh2yi4zjULoti3YcGoyI
oct9qc6XKoJpU+dYmYM/gukbTwvppCFzQvtJ+lx2LO+GcPvd3HLcVSPpzzul+6nHb3YLsSoLzMkP
d17acod3g7wMvFFWLZ8nLId6UYhuFtl/wCzFjMUe4qHszuDp/vQn5dHLS1tm7fxjca8uXjWSXvTa
P1oI/XmopSEPwmV+yXyPTKL6FLZMMX9xCObclAfVmJLpHU9Ry4bxu1THe0R29443U+b0ItnzaHv+
p51bg+uF1Qms9LNGoDepw1zZyO/XZaYNJWh9HT8Dv2yyTzNDVm+muJxn7V6UUJE64vhAdHhZmVd8
XYH1CjeNs9yOy7bqiRarBZlwV8c/hwV19eON5LlCqGzVSrqlPrtGcJCaHA09KXLimJlHp0vZwGN9
h9HklMoE6ZAg+eBqfSlvqyAw52Urooq/fdmRiauOZnXMMCS8REacyVGDItzQHsHbouizNYg5/lKl
ZNCeLLKetXQWzIShsfN5zArWTld5/IpkkeTPWe2LKdhs9kfpz3V6huMvI86fXSDhe+PjOgqYd6La
46dbaWN8o+zt697u4JN/LuDt36blRPBCbQzsaaPisUJuatRsdq+exC6jcTffu7uyTxfiVouWhufZ
PjMDY+I/HpkNLDItt/h9xowVrSphyjZyrs+aqiaL+vav8IQIzbpD9HGKs0m98847ePfherXy8YYG
ZFs5XFnm/aS3O+4enmIRwjxDh2c427Szr9sfV4Jfo/jUJrynSCMcsrtJQLC11WvRsYZg/mtWFB3y
U91yckoad18MIbtRHOTM9/gUbriz7BKB8kAs+m6pBCf5tg8xxKfT2d+va4qbfh9IMUmgCvX3n2IA
PRc6ajYTzrJmnXHOLD04ChFpXwFaHd0UJJSUVr0BEcqoqtmmHQhRE1CB3LXttdq8TKcDnmVMr9Ch
82XVrUA1yEKCzAswUcYJMaWpMJClK7FCI1MfwmHdDCNEK9i60HC2q+tIX3AIOBC1uLbERQaIEtPP
QpYRAen45n83S3yrDX7hINXP2mnTw3pma6TpVPzT3kBVwO2FYckvxumleeSoWRanUK7D2UA0C1qR
69MOYHE6yIqwnWu49Kz6GadcQv4JS+ryVqhwF0FtQp4bEmwmq4hbRu6HQzHDbeNOs06/ukPgywIA
8qJaRbarfuIyVc5rMDoX9uZPzqRhHq4nNwRA1ZlwbeEXU5/RLr0Bi/BgBRg2mK0m8+k4fEMLrHex
yfwfHrFIMYsjdHLckS86mpKRP2TtCgbyLD/Vww0B8WPisT+zL+w2TnXy8RkcN0L1ivpcnhZTv9Rp
WXsAE3z0VBBXdqyXXShdj+YT7KwNfs+G970iWcekdO3A+9Sq8K+B/PujJhknE/g/UCtY4W6pqUCU
dDyMAT420xz6rom935IHrLpSPfqY/CvkUcMcro1HlshzkxLFbJltdfwrVP+i5MbZ7QIdceTzPoU/
vuUoMUZpJL4PUT3m8Lsc2vYxHgD8gfORWn4DdyS+KtVB40SjDhUhHmqAEkH+/mjxTOxC1kqkmrwX
Xzz6LBxLW5ZQTrNlJ9DwJPDsRul32VtiBO0Un+ObK2iL6omtjjJ/VHtwpJDttQLT1nI9ZLLoKSp3
azWA7nRaAkIVR7R1Pjg9dn5ZqMkzUChJ3KZSooiwNzBQv8RA4o59toKS2WiyHQYbjufp90DhF16n
sOYkO22Ssi+Jc8NPNF+z3cz8wr7WxFW1AMVHXyPrNds69FIpFM30MMjsGnWOkjUNGstam1jiOv42
QAknPuQ255kSlA8DfwxBB+RVm2dByYpBMWl0x/yGki8nOj+RA/Ym1L8LHCK3QSfamr64hDy+Vv2X
MLwiKOsQvDOCOAqbS5GLI6KWgdQqdJBST9Vb0FsXsqAAodcrXW/aycaAZt/SelF+u8P2wOzy5qUP
futKYsSVqsdp1YwIj/Ca/5w2qvKFXPLTaxH7o9ukqpAjFkDJUIuwtXbr5vCg43Zu9cJ3W0IdFjnL
ahy8VvRAH7qW6L16M4VhGd8iwDCs/GBhsDMjoImU0qjaKmQh4VMyzyhp87gHWmSfS2G6bA+lC6i9
yC7gX60knmq8ZUvMGnjDOXNVhcSOS0fC9XD9+q0Jjh7lJOZPfehtbDvYL/ikVte4+yhb83ZAy0bt
APJ9qiQ6fzcg+Eaa3QLO2kfncv1izg/sbd+QbtUdenZPD6qI4WC9Ni/UxAwON5ITRXZXubc3OQo1
dsusqnklcL2g2HI3aKnAnBIlo7Cs2HWzCp6bNCLyi3R5Lh6obDtrOF5+FiTQbAZMddBPJRNWQEQv
m4lAsOhJstzsmfE7v8schdIJPmsOEKiP0SxAJNG2Nnj0nReeZJkylM3SbvT/du5julvRliuELqH/
5BYda4pNS+ftJccpu5MVt1fWXi2D7p4PgkR3o8h0PHeBZN3Fsgv1ex7V5PEct/dupbjpCUOABmRX
R1mW9gfTRrz1EUk9gakemTrNvAkXqe++v9RP+TQWrN1Jbsnh+6EwCnYaKKp2ufBq6q0q3aSwcRjk
Vzk3mD6m5X9Y36ZSKzh/LT2vYyH66pnSRXRyJ2KubCb4nI4BBTNNdsYwsX2MVkFXZkoF7KfFMwzK
6avg011CRQ+1A0Ryccr1EogspZpGEwpvZAqfGFuDJrdT84k76NBMxPq4DoLvdyoF8WmtCJmWOYQ/
hM27kRc8q7VG/Ig2P1hUzirAvt0xZi3HCvX81gXwrDXrAMfPQ5x5b3CYDrFegDm3GPayndRqceFV
3JuhNZ7PCEv2aEwLaosdexY0nfT9DhGZzgKg7uHgFP+IStDAIsVxQRLacE2EYea5Uvk1zV/hmiSG
M5mqWR4isj+dHWM7wsaFbVwV8pWYx6UtkoUdUj9YpfRBPi2eac+ml5/8nhLfErbJYRsAb6Estr0V
MC85r9nG/KLgtRL3n6esNgfHVb5pSD/i6KlgewOe/5Dh0nSTisgRD7QyOaVhB3QRRRsM8hxycBtT
lFxIlVLz5P+8Sjwu3YEIapCKAf4Yww6yu7Rh9pTnAcVlctlNKvjUZ/JmvLDF28N/pVe0lTxxglOT
1wkQ8ozcD+KAQ0dhrh3XJzzfAuaBzpPTWvTskwEeLgvvm85wfELBUgwCt2Ti5FOqk7owWOB6Mk4j
Xon19Rf6MqgOVskVrrkw1YpBHLYAYxCQGnqg1TMFYProfP4FloRPNkaDnwxGQfUZUBl5eP3m/a8b
f0+HgjNkjEg+t8R0GxtgrVBHaVW++c6qjxSPCseQvdrSjk8agOg3Mx0WdJHUF0lCJEKv03LNuK0b
X2go9d1yXDtXtwSodbb5szw8Z0R3RwFEQCqPv9orL1QlZ/X7Xz9sGcjZM+iUXtUsIAIx/XtxZm/l
wtcPzarBAdnFN3UPja17n3Iyyup6yEewH3tmJl39grq5v5n0WR8UvbYY3+Hs0o4uhFE3pll17KLM
W6vvfe9pMUOxwPtbHupvZQkBM9m8Y0C2I0p2hyPF5Y+sbkbHC6HtHERbylcYqROGNvqIoxJDaVxO
mMgPtTtaXNBtWggf+whoKZkW1jArGBLv8elYF2kqnsn6QTpC+/ZyFpFtRSJAjlzlgItEceuREsz/
aDzdoS9OBhtdmPMI9sWko8ktahFy2Uzo20gv6AMDMmjki1EJEs4TOQwdinjZiRboa+FpOWKlenpB
BBJH9J2S9GhBgx5xU1JIuldOvcfp1QiP07tvnYz3XvHPEFEKo//llSSYCKIYnX4Dz2sKWah7JJNl
buJ/Ad6kvBreLSVmC52hNPr7/05SotsBoUJ9ItO/ANsqQh65kDf/PB2RUobcKoUsY2HQtTzel7pz
p/Mp0yQrX1fONutqj29AK1VMI5aRNKoH5Gh+JIn+xTuoTjNGgZzk2VGrRI7E9eWzdof9Vs4N6dMF
MOUyzlpNaRBrCjnuqoe/i3VznXk15wqe7j4PYIU9HZoEmCIQvb0ntlfnQcQioMfI7PJ5Et1euoW0
had0NvJ3r+xNCfjooSyeNCvOqWwjineOzugtG0moskRp2bw/P+dcD+vQLK46sbsHJRWP2hZEPQd/
hysZbMjbQFilV0/r0/LGn2dMZKHInXnk3YTWOuNBPIHEvJPEKfloR/6010LuZmCoiF7ZfqdE1ceS
zpEUUftUc1mvuc9IK0XsZ1DVaiRQu05TSHdAdSHMZovrl2UOzAookriL9ZxI0Xh+ua61vtb0CBYc
q0ADIVz8kvwVl0BgyiJd+EQmGbxPHAo3rTc6rgyHt9kk0yKJfov3BYXmZFPlTMr3QLTZ++4KVH7K
w8yZvzRtd/t3V8tBKjI5JoR6ki+NvhafotdLjnjb881EEu6grwYsn71ecQtuHWNVFf3nxwaO+Iv4
I2xbQh8H6Rwq0TKZ0gxz4v2EmSI5Mn51eca5/5DTpjTibFFRV0bQ6W71rWCLhHI0DA+GMumBbMl7
MCLf72eQtfmHF2IZYBM9ry1vB7YMW4NiMSescZtlxdcjrlXgg45k0newZv9kdYRtaKXFXKpPDSiX
gRVoDJJWGsGcWwfuedYAxlzPF/EJhPIhbQItuJrmbdQ6BT/wbNrkdMw18ED9mUMpO8qqBY87jN5d
+8g0y6JS5Tg071U6N34xGV8EuCCCQZGcUaXk7gxcTRpiNRLWyJ6J8xwdmWHqBGk3l8xZVvmk28wX
RBk3N3UPzNEgphf6j6mExJbIezc3/TMFgOymrbAtd89Mk9aaNbdIrttyBoKvPSFoEdd/uR21sSZS
p8EdATDl76QKIGhw9XFCcDgIgquHZ1SL+5nAXT1xdbWg/NcRsqJBoE/DeFyNLOuhdEp/EtrXnVuU
nRHZEqb2G55pWu2csznQhweH53FAgxBPSCKq6PDAV9O5V5hZIVDgFlrtkSoYI2UpS5NDPeGKYo53
dUBghSDrLN0BGPIl6rYCHO1AhuElMeEB+lAxcGbd8sc+uNF8II1GwMTW2O7rFivVOU06inrIb2jL
mV7bK841XFgn9ccA/QoIagR+G498xvXaPYOeZLYW9RI11eJz2neMx22eNa5VWkFnstzeF4JLAeUc
EunlVvS23GQZ1Di9n6Rh2MWiQ1WQk/owYlLRQwohknDBet22co8u0P42Kw+Bi8M7cHdnzrt6v9Hd
NaLxv7qrG2Ndnf4aC0jtNGPDB6iv3KKOPDRqJmqN/CSjaME6ApHUhu7uC+2devRNzleGcoBT0HRp
xY5JEHzTq53K/fOYYjzrqexegL8mAs9n+aGGU4Syg0t2/PYOJxml9Yir8+R6dIKzfBrYONwiLjtD
yFDqb+ip4/DfYWcWO+j2eZTe52byTGk11tWBdFNaMKi7eOJ9tz31oxtxAtXLKA2wcxCCGpY4M6L1
TSVA1WX1fuZhnVH/hw7zQLyey8qr/YfG6jAhdK1aca0HPX49D+/E5fU7GCA3s5rqyke7Z8km9p12
J4EcIBUtri0Zi72CtSx5BXT/uj28WkuHPn/LOX1TtqoFQGnfdsBAmiZykvyEFj//14X2Ohi80LIF
LsK9woBdh0bIFiIirHs6io37tFQVz0xGh1ZYdV6KArftztFtanScAptyjlmVSnLodM8/ZrbAyqWr
4IOPkGtdRT5blfGXnWtOvmbgzHo75U89fTGVrxqvc8kom7svA4SRkf+EVVBp4Ej0RwE4h0xZ5JUH
yyWvQBCF8a6egfZnEe9kEPiKjIgLuADV4E6eOWZScq28e9QbtBhNd2+ikpGd8ymJsrLNJZw2wNIi
EbO8FZ5vplfqkcoJSYzbdLgyfcGMTfj7x51m7a4BXDfcpwtpcRS9EjEdj40gzLD+9AXuQPY9qRia
Rk3oFUYQuMdRVHePhfh9ds5nHiPqNjnCIzfAXqrepaYHE9x24+ZjdkcxUhejfYVfSrld0+ecnIDz
tGm47iaQCHy2djPXPZD4p8ZvWK2kskOK0v++3iIMxoPURgLvpnSj0MkHSZ7HJzd87F2SJoiVuED9
eI0p1gz+Pao8zdCAejmluXoThp5cIVgKg4Yc8JQuxdWiVf+S8NAu2lmRk/psyVCDnmZVwfDhrCxN
3z09GK1DdgaTeHvcOC6mR9gKoJq5+bQE2WEhKD6VbSoS0tMwMKRLc7FYkg91tO2E/LuHxAE2Odgh
Dybj/W9v/OZBWAfhcaR7oc1J3I5QMJFyiWFQMlvIZaTXw4uzblUVIi4f0DFPYUYScIloKcNE8VV/
8Fm8kEfp0/2/tB370j/2a9a6p1xWKfpzZi4FEghjGmtxeC300ukzClwl4uFFvhxpzdIAyPByM9IY
siqPntJeLRnWHtD1xRTBBB4yBa5e1mGWkELkw+OjWORZALDuxahKgc7sIUQtEpKpww81PPHY1WZW
Ke+8JFHIJD5HRX344yNE3FdxsxKYA+4HTmZ9Gz3WD6gXPGq1Ht0c6oFa/gZILgIKnjP0IMHLkwJu
dgYkWP7Ae5VUb2alUowrFhHoxIzMEhase3d5tB21mONRXbODvxNoKaFO94RNFvn+egrlNkUjjI/u
TjbqQYuhacBbLu7CU/tUhmGPCbuDpqcez53gpf3FyeZJYORSXTjyl1Io2hWFYAJCnrxpUMwt7XM9
1wbi6aLi2oddpI0ARy8pqa+9dgu+5ctNfIH/cizd18u2obSgaYnaBwRX8SkPASEi1mdnCEerizx6
ASyF/rfNT6sq9dpHdQc50ohxc6d3xkF4C2QbzNRpjjZ5UekeUwPTAKGz6qr+igP6TPYPVeOugUwm
aLNPvmvErHE3scfyWgAotdHqZpJ7BA6RRDiQ5ALL6IN65H9YUdrZWu0F6nzOwuh3uNRqGVVBOCjg
A4WAStWTvDGLqwVIktJXH6cevgeT9q63oFis4C/cSps95wATka2HQPXVVEa7PIUv2ZzR3c9g3t2H
iYB7f2obR4UJj2fvCTuH8mVMkrfyTRgXYDqleTGFyN0gxl0TFeM+WLbpUL2KK8uJfUDekj/6FOw/
By6mm8DpVUdLmK6qUF1dd3Hef46vZbZzfp5dRQ0xaaPOtydQXD12TxKFuF/gVyx7gYAxvaHUb3lu
sGtowcSiLnt+7Y9SLJa/VxlfilXypnU6Ikqd4jDDZVdw4jMGX63VsYfFD/Nqp3sUQj3o0ZnK+aaB
xJnzAz46S4wXApUvYoc9XAq420Uhy30JYwpMlEDJ2fhqZeMhejpUqxzv7h6M12SIgpmLH2HQsCy3
nc8nn/Mc8/XFi/OKtU21vQgRnvSNLeiTEzPx18nz1YGX8+ivjDx59qTYZbjCLWQ/iStL172iLKAY
MTZTIVaYy2joD0uCJtF1lM8N7/wvU/qM9nDkvAc+Rl5j0djRKAFqintM04MJkmnGCxOuDexxszyk
jWxRT5JL1uJy1IyO02RwlJ4kdKSyAzZvIXznCCyzUtyE4pKtTIduHxb/mlpBuVGn1zPvHBhEJsKW
8z1bidvvIxc0pgkE545dXSfMZt48Nob2JH7SlqSgt2KsJCwCGxc67QgrTcxbhkTarHiaOFZTMuLp
L2UZdR1dguR+m5ASmy5gpkdEAvcyw73aacko+spL9rMRIR3RlpKYAmHXXfk5/zpRHNvtIKM8IVnQ
11dpko/o31C5VYiKHeuUKKmhIF6+Ps28UZMUGcXg91eMv4SfeoplMKztij2UTpH+C5G9DaODsEtW
/J8Ar5OTAmudK6+AKaGfXl2Gu0SnXAD67v5AfGT1IkASEF4Is4c5viJLdPic2H/yvzm9UbEqn1j8
AQi4X+HJVlBB/3Dbduc8DUFQAgc5hVXX2XjpTOevF/mLWcTi95lLZ24y/4Y3osVUJ6bE1K/UW6PH
XABNTPBI/JLx/6FEv2WwzAugGdxo8+rrqAb4y7vC/1EVm4LnmZah3omqM0skQYFM9mxW071bNaSS
cwE5TBeKn6ZMQy2j+W1iOpB93XeiA4H2ju5SR1yjTXLyEegCEcD8VP0K8KIqYZy8fubZ5tRZk2KV
SXTSAdgH8P7A2FbTn7ay6lShHbxwT5aSm+JvDW/Ur7+ZSEC1lf09HRX5m0kkNiydyTRaQ9IFvNqi
tDX0VoiRSNYyl0UIOus6f1k1kVzAVJHizEPpyB1eMuCduv45cXYdGnIAeDpWemUfuslYLWAFNN/T
yKEI0mGlw5DNCberouluqjddyPR9pzkxpZsIRJG3sy2EeqBmwNCEt3edjvA6FYoXq7FN6Bc7Tze6
f+21iCgajAc/YD16iao0NfLwvKhy/+UuOOGPM4HOszfSdPRPRW6OZJOLsFmUh3i0A07k0vU575IU
h8mHU5LTObAtfuzro1JzbYWUSpkvMbqmdDUIH7GFSR7UYGBcDn11kxdnzlxPBBNcC4AiJ72dcJ26
NU/bl8uV9T97HnXnZbyiQsC/efLppnCwrCAF8cL6fGOaoAtVB7L8hdcphTifsgaZtX+detiz6rQI
/6bxvQzt3VoIxLy00ma98gvn0BRhfSXAaFv4iD5Gos1bJ4JmUwfmooZVu48mH8e9DUMNbTsX6HPd
wJdqpQVmf4urLGemCFaSmk5S98vVk4w+UncOXoE/RezpZGMrWyOFOsCjiIokCwdt1gJSJstd9IqF
YcJG6MNGEDXjlrAs6URyV83hK4UfTRDXovnNsZE3Qinx/wJMp/JiMjxYsQWGzv7kLErTvrLApYy2
toCpoAZoAnk1koXzQ/8JxGgklBV9bvQCefdZiMqj2fpicowtt/pl/Sz3ABM422WrvPnJBnOxwGB/
yNL26cGA5wSR2aWgPmVteyqn0L3i+wCx33GRv5lcmdTvoADYqroacLhIyvBSnR8ENU5vTm5gIA65
hJj87BCGHquhcZI+MZI/lJ9oWrlLg8uPTMPgMb19hzP25Of3TTG8ALpRDTgpnLzNFHauq5LB/Acr
4xlxahUxmG8rxjELEhZCvXNkrDaOaOle6uqe3piwkf8ectY1v1kbAio4+znZnuW1YvWDBilArpaD
3PanA9VSoIJL93MIB5Z5cSEtiOdG43xu7SdO9AKoW20qY3FByLh0ly47lp5tvrQH9emt9XMF+YKM
YE1XQgTuI596WU4D3d06TSTvAC7RleRsF9Cm+k5e36AkRJdJDWShPxHg6t9VhOqyC6rE2P0izMb8
GrkuEtEJ4GRZH0AILDewLRofATV/v9gSxA+NvBglPze5edN1SQQ9FmL5Gxky7xHmCd/9BLaQW7b/
w4lx7nvq1HV4FxVfUUrTgJro5R7sfqlFUyc/VTfsZWBMnNdeeZH2Npvud0VrmdaWggYpsX940K3x
4GFI99Dk0/P3r/BtKCXnJw2TKLs/E9AFo1UoFCgyh5q+GIFn4zU604KklRHMz0leNBHtOcYpy5Vt
C4AfmS0sDlGDqaE6+4yBuXWpiURbxaU8UtpH745Id6TmFfz197mzaePnIMhR/1OuoRoiRw+qITzd
5bm1MYDtJ/TPNAuo3ApHLz6uITdOOMDh0eXzEpFnMczyzA97oTLZbKuYPr6qR66H5YbyXg8WExUq
TeuUjYdiv8986MuAqctSUxJ8DmjPNwxjh6nYuGVDLxXM12SXcRkpWkp1EtT2LSkfAWO8lEGVBsUm
O19Xa6i9nhUm61Iu3KiTC2dM4OIuX1QGk1EUPIwdYjapI0IEikkdbgAlbrZH4SxkzfM7UO/2QpUX
X8k3IAzyn2dQQ3rLbX1d0iTrY+GSoGJiBYqdw576LWYCfmWycEjV5yzj0clC48qWUalGGorDHNYi
IQIe9w19gecJ+xFDZim1RqGhSAjkg/Xd5vBmNRRX950uJ7LR9Lvk/1p6M5qmkvY9lEnBmZCWibLm
N26ECKyeb91ok6t2euzgZ5EMiSNGt8DnDi4F/op2JI8AbNuXQBuNU+/BbJcZL6ufXU73vcDr/wfB
omFnuU8RcZ7BOm+aO6jLqUbxyfct9asCTh2XFmotWqbvAHZ4aq/iWO2J4aNXNaes3XOXdl43fE3D
Ysljj8a0at7mKbv5tKRj6xdOo7FRxloq2eonY+a0WV6+2ihMixHEp52C9Agk/osy413o4xngA63F
IwehpcCW/jqbqmFRrfCM8fRq0TV96RSuZxFSvX6aFWmD7GW+sVmV/nSoOzO0zG27TSNDBTL3uubE
yXFPhHuUHVDtbUb15+fb4wwzk5m3+Q6iXpRChbhoQYvblSUQiNVOT+S5L0XIl0et/BDQk3KWrAs4
3ZHnapycC+vap+86Ve2J6YG3pZ9h7ogYyg0WJx7m7MeevQALUubGExO7ZXqaXT7Umfo0pagfZx6c
GlcjJQuy5QWtS8L0+fMi3nqTsLVml6M8gzEkMU9i2mlxUbxJezu1eaz7JK7b3LbBuNBBITwp6tWe
wNyHNhro2BIruyBdtzpcfgtfxrn8lP0mA+MMkM/7Y8IRwjVio30lf1DQhml+7Fnl5mw7r6gB5yqN
sWcUxT6o34/sl08/8IFdSDjDmd6KmnTpuAXQkgQINmH4YLvLRVfLFmWWDQ3icLlNVRkXIiWk4Pg0
tGOANNUuPU6bcPcW2Ay+3ZNY6MXPU0QNf982sFks2zN/vxAJ7/m83QaBgaSrqUCX5GAWh7u98cIB
BS+JSjMUELFCOtJhWoGafE5rrrdlZkZZhffFAXfpGi/WkYNgYGXG16J0FXp/+tDnPvB6WVQPT9KE
iPdhYxWGEnJj9i+QKIaFYnZ9b1p08GTvKPhzxRX5zqQB7IiNa8nBEqHLEwYT+Bk3rznV2Yih3zzN
CozsI7ZtSaqkJFo3a5BnJMhtGVJ1skA3NdPlJiwiEiYFABfYLpabb0ZkgHx0/KbGUZ+b6BnkW9nh
IKSSmW4PMkDCVeQLhSiILbdH7J/5sL0ZZXpVuFedhGIR1/XFH80opXdwYFaZ6UAL+DUV/BPnFwXe
BFlqRempAzTfCggee1+gpJyEK7SpeZWiWlmtMsqlrWX5fsNiLtXfjFxiT7uPhNh3k4oNGwL+e5wD
akohSeiU2p4B5MUtXloyXcSuZSEymr6JXEArWGTc+//bWelpn2ePoPz4qibKi47IduZ2yMAYCaii
0IK65CM19xdGIvD4sVzCFBU12zxM/xXJZJLLhn6ukIO9JoLpqVjVlhvaApNWRRItIKS9It4EJ8yc
Qf5BA9TuKpTfa+XTms1PEYmQGEltVoCkBPIFv5nW5wrEcnyZiWh6nI89B6b/14eYvYalgCCOLkle
0jiQ0RtPhSpPXQSLqsscYo9eCc2PzS50LhpL3XjIkLyVcVPal2qu8oWbMxUNjd1gbborgmzMtqhG
wGLALgcFCHGeRxIxmlLlnJD8W32mv8rgf7RMB7/jyU8N329e/O5N1s1WhTXPpBYMQcUEQrgzTAyT
BF7l+IhqobzVtyEokaKx/TlbZJAjyFqSUnj+t+vRlg7yzr8UxTspBS7dbJrSU7rtgsFdqkf7x0X/
sP3eg8GyNYXehlb3f3i7366Wjy9ZBKfuu9omL0k/9i/CS7kIPacBmgE0EEUO/Udo2K6Xi98CNpem
tckIOEsGgalDwcHDw8PizKpHk04pJyYn0x5d5sFji12Pz49YCuKsgUzfo0ELKEI5i5Khm2smZYDB
QrC0qzhDUM8W9z7IxiK8IQNQiXOjOhwiBspenDI5RnBv5frzXrnbkIJ8CSL6NW220mESmAcnjPeg
itn+Nc1dXR0Djt2eIYHSJcPZtycCYjUhs+uYzd82kmgvb+/v/wx1xQFfixDznIjHqOOO4YEEd9O+
FYA81V6gC4Qbq6VZcGkRSZpDZahPZf/NhhH0eLRCmwk/Z43X+mGuU2Y75SH0GNhJXB1oscH9Y4Cz
HKYqtgb74Rk7nIA/QdoHzQ/W1kNVl31c18N7LoAvZukXDB3loQlRGBphexf7Z8q3QL8ZjfwpIj6J
tecF8Z+b6BXhJ0c8bPBz1PAvX5LEHGOtYpp0mRFUKRcMVTGd/sL93pss0c+nZI8+w7s4jXOHhAWw
Cvr+00Qki9HUjtYqVyrs2PnjnlC6cL74HlcmrpQAG0ENCgWF1I80DmtKUfs9EpaSGAg24vzI0X9W
c7olrWHfEGmmBIk14+HFWAsuhWywE3Zzhz9+dtnPZsrfAXAHDugVFmWB+zLo/u8fl0h8B6AhQrma
gIafY+ugh4uUkbSZsFtWkfl30ptUz8COA1zqzzz9s0FqBCDLfNJJ9A8QafDpks89WGvTMWbdVGr4
lXjyhkQhzBr28MKYVQQOZC42Ytz4CQCdC0NAHv4jOIYtlIkTPVfos7hf3u1w0rDgel6bZx/jSaqv
B/oAFLlcBvhSgs0foavLXMKx15SWZwAGcc4bFThXvnAFeSNjqnax00a+F9vzSH7UGMG9WHsHqTGy
fj6lFiWq3T4mGbOHygVAbiATeUYNwnPMLyQzTQ6v58IB6+6PEGKTXJkn6uD+bqQBaicwprmPSr+N
2xvda2sJC0l4WIdUK6Quh2TIMq30HNYglnUJhETKdzWjnKcj7u0nP2FybfugCCTEr6YuSMoD5Qgu
fBfmBNdRQOpolJjzVFWDKZbvMI/r/dz1f4BxiTkQfnfHRApe7y/8D4+8OwVvKqD0Go5N0L7ZDwLj
fx0izI1e6sLwB+9mvEszaAitvl2GcFhoQgJGkY9+B/SKuIAV42RhY9PQh3fRkQCkm4Ei8j5jpIPI
vtajtrGHUHBfN9gJf48keOt6TeWS4u7e54hSfgE6oNgNBfxBlpTLgkx91GbzL31Yl6NkG9t4Zb5f
V2gnia8bCPnPJAzi8r8g9Kb7CE3OlFdeq7pavUEd/sBfQpvy8rYNXB3p+Mr6xi9Y4cwzITQosd89
Jekjna5BgtyjH1Q77//UbYbS0jXdjwuN1SiihNq1MQCTantA5ounMoNJuVHsl36/nvTxulR+wnmi
5/2OqpE8v01+m6e9yI43r6w+RdLXpyJTNB9+Gm1Wwb+H17T3DTGHBUDpUOPuR1LTD+iOxZ4d7fpH
rQSH1bU7bHZrXhxnw4qKNZvE1u+cc3B6YUl/xJ/VLh5flewa7WvhSszaFFw2MwX1gCAMR0j87ZEI
/jm5mSOuuHxrlHCa+Wn23conxqILoF7bE1sz2lQBxiMqEgRRMtQUEZzQTQrlBRSc6ru2Oo/UfP5j
IXbJTiwSGG+GQKz+D6q22tJP5ubOvNGYJ9TKt4fPGICr+ZrubwgMAw40F6sz9UDX7fSvv4kXAzDN
2oaziAd5msbhNTsD1AqkAbD+WgtQFJWLG+iinobguOvqjKTtxafMBzXgr0qy/nNYksnNkF8cO7Ex
iJL5DP317q4XREyujoxHGCxbJYOpsbxJ4iO7LAbz+L41P1G+BYqvLQfHgntQWMWY0xjClEdA5V0c
wrvJWqc+FxoE/ZqO1RSn1DP9OL/WV0dVh6Usx2YMrD9xYvW6Nb0Ju+xqEiU6iO52kJvX2zoNt52O
fL+Qgd1OA92tcsA+ljeBiO3k2RHSHzvFUOR22RZ0kRY1nTKupYQth5wDKsNxf1gqXu+RGe5KXLPb
oe1zn0nvfd5+iUqrtixrHrgi0SvaHRMJpMDc4YdVMmVjOKFgj1sLpo+wPvtf+8v/GK5cm2+pCWqA
1ExJGhGDrTj1gIJx/sDtC1QhKuWE4OQrOM1uQfhOlNj+GcRI72jzs8qMKx1rE1FH5kYEkuY9REHw
5yAXqAkxTYX7JSnPHg9qXDuP+QrL8qfcRQyXbGCdPcpe0Qfq7FcR4rv963exdyqPDF11aJW9rhKJ
0zQKf84Jg4ndzpGN8bXBR2uOhD23IybQL9FRTteL5P0uSDHXGG0bVTs4GboRgvVuiLSLVDqeqfQS
KMwbBaZV3bCpfhaeySn6D9INvPI444Znty/XHAK/QNXPYkrC1uE/LueFTErVQ6+45WljMU4/PGN9
a/rL/CCuQd1FOy5UFmXdxptxe57g+ImMM20tK8pv4E24/CExJHz8FBuKvwNcNYc5/KOHojyDFP3K
wPxl2XII6z+LHEGDfdpvBBde2//zswgXT7CcGlCvTrfFSwEcPQvM4VXnziEjyN8RoRu6DTA/mNY0
m8EZudeW08Kq4551bDNshlKmv23qaNodHE0SaVyhsKKF7/KiZhbGHSd6IyTI3xOCU8gEzegHyrSp
Xr0KKH3A0ThxFm1WOLEcTbbxL5OCX9yBpfbL2ykJCJZNyiYnbbXZ0eDYjGkVUAjCIktPhMFV+7DY
WTGabUqmzEK5yiKavXEasskdtUWeoZRoTXn5SOR7vtWQ5d0MQBW7+Rd64eVlo4THrC/nrYOClzKU
lpKquuIS4/OU/GtvrzWOcYNqPeguj4wGxLot2hv9HC3KqwdG8PDEfqrzApHgaoNkFY7QYqnvMT9h
4NC72v4nZYWfxLkRlpfTNXXOQvWJyt353KokQcwIQ0fFzhcgFdAHeW2wmdKTDo8BW92BoKSD2mMv
Xz8ZIj/RiiOWALNBp3ZxH9NM2Z4ghPxxrBrj4UhpiHzkVU9mMSrNs/T/VJoZps6HrKK7i5SkLq6Z
SYp9QD05jirE+XEpKkZuPmT1+YuGS3smSoEOj6SbG1v45PD+XRO2vxEQCClYSCVe4WtiQUoeGl2D
x/8Z6PGIwYjYzAPdgCMa1mveTpNpGJ0HWy+KI2L5tuL+d1ofESgUq6m4XigM6uS1Qy4NZOnHaAwT
oFqJ6BeRs2MoFyjz6f1+8hvDuUnzlBeFljIM+0GnLYvDWEIF193S+Dl94XH/GOyy0N1v2gb7/H8P
k44cqgYvQXB8+oWBwsx4OUkN5OtWKGITwp1f6nia+T1eJr1HfA5HfZkQnrKHdmnT38INKlFB400Y
gNz+eKTBZRo9x+NEtjEaYc6ULUhoBO1yK810+QJCcgwuM/GJfvTuWfka3pkyFpPRHZN5YQT5gJ7E
dkCFoD9fmR2fqXElRkdIVRbj9vqbRVd6buY1ZRvtFBK9X1OMlvtE1MsWMJYE6KgpN/Ex85RMdyK6
cUztmaGNdHCC7sjlQKkg6DjjoTf8wc80EWtVYVAtyNGfCjY09JEm4AGAvOgvNqHuZjO0TtM03BRU
OrmtEnk/JjMK29E/W5CWvg9aWeGMLG6cig9Ci1cRCLZOhj1OfzhGLmqC1AI1jRKUQc6DoVfiDHPG
HD6HbuF1Lp7Fr9dl5m8dIWktQZ5PzRR5MrD7u2U6To1vYeTN5v9OceR0gFIcNccLM+qF4kM2AjOl
RB8Off0O0Pdynnwfk6KA+1rQuopp72l0wOB6wjGoppC9RCfCcIVKvHd0SH8tSds3lITzeD1Ax+XQ
GJGAboW43z0y/jYrFVaK7/HGs9eN7pRJftJXtwESld7bZ9oRTaJx2pSK29Bj8cPsWInWoc1LqdxT
AnBs34EN5d54h2gOIf4hYVRtq7IwycPMUTdbTD4yPG9Ma88tlqUyjtWOHeGSc9EV0QFd0AFwTE2c
j++3J6N8zwymp081Az0mO4FHaeflhwf7EWzFUEkZwOiDW53UlG3gMAxSUDbWpdztMO2/8SZ3x/Q1
FPy7o9fIi57N7gsT3q8Px1nKHgYK+IUSnXc9yiTmv0wFltYF9rm8I/5zCEpk5WypiBIWEUKNjrQe
ve6mX+f/ntKH8soSUEFavl4i06yR5cbWdUoQviOeUd7iTLOE5xfwnY1vQddLsvoKanBvuO+uqv4q
T3tbPZ/KUO4GLfsMg952uzxSYrukrG0A9ORAgzKhT/wXZDwZWf5ULyZA6mn8VaVYqNA5LOACv20B
fEOJDxT780h+NNccc4WGkZvHFub5vJOrjflAsABS39E0QOyPvO0JFgadlN9MRtJ0Bl1Vk16X3CHe
Zn4G64fhuhD/v67A0NjXNWqlS2y6l9KuOMj8DxaVERGFzPeTnowPq+c7l7ALABD0xlwmXiExA9xT
RPAS2zHvwHHkOREXbVeq9bizL9hK8gTcD1Uk5Y6ViFaKCZn3SkHIaYSaNQKkM1QgRtZIiaE5SxAN
50N1wAGkhPpSdQ4WVU28crJlM2DK9SXqPtXyF1QbJm4Pw4vd1wK2ZAtL2N8BeYD8htp3DLcxzsKj
rkbHoTYuVvQA1Fif+tMNzFatscX1/RYABChzTjZareRprwoQn8+1gwI6s9Ae4+Cs73+g5Uswt60s
6Mid7Aapsge8U6T1hczn3qrYQo8UupfMdoLXodb7/JMnVbgEZGx9iOLYVE6e4rKsmwVMqGk69agJ
1UcwyrhsT6QxeU10bKC7vwrhhhu1im3PA7liBljeX1OyMhBRFy5EEC0pTMPRCTM4gLlerL2maowI
CeDAH15COhgiNRu+xg9E/qqgOn6A5uJmjZTEnuiuEECeH06L9l4www5SakVhbz+Y/QanXs5a9NsX
r44LNx99mvbee2ogP5uQt6pGQcSADDTFPGF2zTMeLj3MApdsFFHTP5XaPMQujBhFxWgpAkb3K0vF
6icWT8+0HicX8PKbgpRyRxG7pwbki+psWTfMvk1YFrwUZuP5MUEuMnatrcguFbs1iZYxWlQk3c5r
x7bzluo5FF2p8HaJ5hsl2EOtzBEUW0IZrDz94KiLp4eE34/KSLXsuNeoI7aJ3ahDd4hNQvP5lWcD
tYaC7kmksOdbeqafh1K99oi/iVCY08liH5pKSctS4Z6/wxFzCXq3VF9VoHWdGJ7crOqNXhtfDNer
dbkuRUvBnGtgldAA+Zj4VMQwhe4oa8aopQUyoJQWEdeRNTPCjbKIG9k/blOpo13gPPZIu/uI6EnI
NtaUiKDS8kHA5W3hLy7BgKZqswv4MdGmJPrD0iGQdzqJfDiJxEJTgxOE4PgIrgWbd1pItCcSYpgP
YLbnmqI+5Rr9j1ByS5PGcdjhk9BmpIzF5pLU6NMjMC21d7rRQUIPma4wVDY6/bjfIow5vrQn65fO
cfCseiIlG5gYYOicScZ2QCB7lgV2PyzlrlLYBIcWRL8E2SZ/uYUFY6sY5Qr1ASjIVnh41z0XUlhu
+cGBLnkDdUtgicZRznl+wvH1/qJ/c4ZQq6SOvSto/JUH5Aa5eY2uk+Pr9IF6reEQhHeHelfmr9/F
5aPCS26iEMZw7sFY9aQdMeYny74w05myxhhIB0WFHhwvXTmZ4EOCJu67S04mFKkNWlZi0sMcFFje
+9DX5gBtZuua5siF4YVcGWvbIQpG8d7aFhG3Z2HaQ3VCWARzAPp70MEKbWctwuXQApu49u7/Sog4
CsXkdFB3jpzXe1LsuhJAtHUFaXPHSbIJ9T9nqOS/aFmGyMedbozRZDuRcrkDKViJTtWolUzF4d1v
IVbdY+jes6vg2Vkfh2+iU0XjYj17vWPOyNCTyt9eLL1md5ic4dkAuGFHXMt0FMyVPMJnBwHEwJ9b
egNllin9w6YjbegUxIRiKpEXQYA+5/N2igVUVT1k9OyMo9urdPDfSOZX0U2go4kVXKrnHLykO487
BVaYIIwCnO22i0zk0lZfBq9gciYoeYhYnhm4qu3Fn3W0Lkcp9w9ldIBpgZ+NA1e77YCaQA3kDGRU
Qa4L77HIcD2QSB0+oIgHRkZ4J+zopPAB6a6aLKqYpmvF9vdAk8YummeODFSTbayhdQMY9wuHRuzk
6roLCnb/Hmj+cNtymrsvJDrrIuZ9yTTy6o3UO6TV9tioybA1kviel9D1zE5AxOlzwRaTtsGH67k9
7uzljWOTLZ+7iAo0VONf+I9HiWwspcSjVcrpdckQVrP7LuitXott3oU00CynoWxFD95LHzhbg+r0
gu8Ytp0/vVwN7Ifej/uTsJwEg/pBB951lYoKisNSYsggpJKHKIvYE6xipxPx+IDrAJ7N0p4yVezv
SGpT55BND+PwFSsYqtjBkp4s8FOJ6DxCoyGiFFvhyPJxfupelKxybs7Mht6pw0m5zue8q0+G6v4O
+RzbXgEMbxTWk6Cw7YwD+10QAO48qHJnSpUZwtvlEtDNrFmIIetSpOnUNBtBS6zEgjkmvdfMtKD9
frDd1ADB7EzSfpkm/Tw6j3+8cKqbLfmj6vD2BxSF+U1PrUEd4GA5wFEJ54UwBT9cvFL9yl/AoxJ9
rUfCkeGR4RhjAFW4T9LdPsnFoFch4uttrYgxUeElulasriSxLQ19AzwNSMWGrJe2SlKKKtuJZ4bE
kKRdwcOFVhSlbCqlIwoZzX3dKDUeoZSgkPDhr+FCPKn9S/o+T+/gSxi8UDUiBAM63iiT+MaVYzyU
nRihrKzy/+nU7LIxoX9Krg7d52yTN/KeGpHUT8zzqWLBGVntURrXL5bZWtQ30mwMBctr7+DIGQrc
rVFGpdP8mE2K6wCrN0EFXQik4pnQ5lc8u6WB2pRlpJZkD5Gxn1wYmHUS2DgMIfld6H2wp9adD2ub
H11mbDyKFE3N9SXSCsIriFClVfvkrEzHZ5GdyA9l/CUHRA1o7SHTzC4O0OjQWtJ0mf+NtQvWAHuY
laljcVdqV/WjXfnE9YqbS9Xi8x8Iw739bPhprUxOCdyC8vMsKrHNDtO3msXj27Tw01Da0bKe7txc
vFWV8e3rDlr6k8orr2u+QQSOdlsF7I00icduENr1cHkAd64K1TOwUtPfvUbJ+3/XJbkI5vH1P6Vz
qbRqwdYqLgzfjBVFSIQpUnIaPhQWVYBolt5K/OQAnjy+pHVEAbaDdx8CsOLoXz0i4ls7bawukLWX
5B8ayNfWlYJLJdvnMivyzTKb6D0docncjiGl6kl4RVOgpslMYbH4OAVmiaYPVb/q5/vfpzjX5P3J
QLPoT2LuUzWTBtiQV+aY/6Ogg/Z02lRnlz/EazHlSK9QsTqOwrXqYSlRN9mPhe0jjrhct71kRNqB
JAvvXXhjmyPo4KPTA21xYgD4xMRbOhRkKG6NDjYybwA/tseQwDKo9vZHonzQ+lHfvo275v1vQkDf
ld73kzKS4dcmxi2ZEC/Uqhf3CTQ7jgxgg4Vt7qTFP/PLzIuq8bEEr+TN1kIwo+6ZTTsJWxPDWgr3
3gb9KDFIpaRQngVKL7zSNrwNnXRG8bfMwEvwFraV85sLHQ90jGivtj23tRwL63w0lDL08kekWPNi
uI9f9O91PRf77q2pVuqGP4IO3VLWbtucrk78GZ1ZM3anVGcgCxeAuidNv5cl39b33qcPebhVrOmM
FS4TxfikBvxMw+Y/3DoIUXfzCU90GngQoYxtGf23hTQfJ2TPmatbp8BBMDmzdCYpIPvHQr3dW+4n
ksxGHp4wV/w8G6FMZisKHaPrKaXPPb39OqaIv0CHDQC4scg44tYBUzGMdI3WJYpXpWgaqhKApS9f
E6nWUag/dGp/qRk6GZdOOmGqXeisqSn5t/Uz/Pu0Ltr1rcj6Q3+rhUSvVr0v+0+CK2ZAYnmaUGpF
DsOczjE2yWnb/4z79j/WerqYs+xOsQXlRApuQyF/0//Ao7uX8/+DhFriUwAXtzjwVM3gwssEfPD7
tZDJz8Y6jmBt9gQ0EXfIezhiX8R038dKtU93kfnaOsq22+jXdB+X7ST5/K/JG19MSzBdK9GwNSKi
/2hiIzjCFrx16lZnKMEw9nCtj0nBmPzn9Bqp8Bjpc2rLWTjRzVjbgibRg7RPR94J4d3o9O6b64pa
kbkVeIA0oFk2dWmPW40IYtPPUtr1y2Nod7rTdOyR8uOJR0qticOl66j7s1aIQI4fxevmOb1v07Xf
FiQCD2n40P9WIgKlgOrstDm7zHb3bYQDZC8Kpd+Fu8DNBzTGG4IQ0Ng0GfAV8HXLVvPJGK++6zZy
bQxetOpddRHZYEVi8JSJ2FepqpRLdxyakOFre+Z6x19KOwp2xHbTuqiI/xSK43Wma2ewDIpT4bIJ
W8wEAqRHW7m560p0qGwH134awW4SrRwyF2lTVx6Eu6Bs0mSfbbycHDcQhBHBLlyMpGRBGQCng01g
tdWzrzYhVZjRnSf2KVfCTquAb9atkTc38aXv+D3yInCL/SXfD363gP8JfAqWB2X26C332vCwigpu
Y8AlZtmL3U6F8l/B85G/4PVTMCJTPtzZVdkfDl1plT24lIoeEWA61EZvvnlTiGH729CeTn+g3n4W
uU2PYxLcQ35lAGuFzkwyuSvU30wo23jXhNKsSZxDJ1oWss+NlW3HUbkFNELOH0wAb15s3BaXo93U
Nn4RdLTMUQvAEfiRLiLf96n1rIYgC6tCmYIrJeUmAHLSFkFVtr0EcnNdf7jdRycFaE0L0Jqq61Rz
7a6o0B9XgZ/sFhS31Uiga2y8DLbbnTk7h5nGzlAblL5F+1ZDL8v4JEPbGJzSqV0+a8WWxb5Ga/bj
s050Bp7fhf3Svq7ydwsGOukoMG/Fbv8lGqaIMmJrVN5qDNZO+Dtxw0RbZDc7hPlIhN5n8o95W+Cu
DNFQOA++SkKodgCIBR5ScPqTnkbcCpPX/tjdveU12bJDD5TlIO1BCrIrChbkKF71n9Ry3m3fi1Fs
CrebDuIUBE+cuLlpZlJM8JOrpWno3qYDgwFttGCZPNyW1yzEuYRRM7Q+zCjauWAQy7t65rP5+OZh
7r/dI8nHzusy7qXBlV+jD4w39tvtCrd1Dvkw/1aWoerkfE7svL99yQDSBr/rkp45tx1BsnD7PQnE
YqN7YVI2jpyBNTx2g4yrl6jr3uRDADruzGkJeKyemGeVinTaxWJJsPkMR6V20IZCS2zJZeGxGVR/
AsPJALY/koCXhE+rwgjLJmqKhzdX/H16AxYcaEBYIsQLd1jXou5GEFRZ+vK33YALwbM25s/9ZqNB
VflEyFPUwkhG2vl3dNo6ku7xn2Rjh9cb7ppCFHlLsog8MdU8/YohTs3Jreeg0QL+B3c27qFS1bnf
HgTqg3qnf+X5up/NBlCL8S2uod1FBMLIXTBgj2FssSq3rpoez4LQVhptaf3uLLLm2RRGuND6maJM
RRICxTe5tn6nB72Iu/5nGaEUtTNmu66ME8UAJK4vaNo7bZsh4g4RCcTjh8LC8C9MAJUvgUxB/AH6
+8OgWTdvV2RQAOcgcOxYXDcs/HFCw7qlECqarKSAGvZg1I/9yehaRX3l3d/ozPgWzWeg6Xyk1ej4
pFA3bPU9vCuHHF6K+SIpAm2pyfA06xQSxt9czR37/bJRe6MxMTMBgpK8u+tiACfAcnLmtLyFQEBh
5wzMgHcxUkXkCNMzzDBqDyofTDIw8aEuPKDanUAMlLdoPKxkOgxDcveSd6QIWxmLXPx1V2AiobRD
9hlqjqB9LjgMl1R85FQ7WKfifnQ4Ws5X97Gi3oFo7TiJ+1j4C7Bc4OOj+88Zy5e3paYTtveQCk5a
YCIztkVvFzmOlaN7bAqknKPP36sSZXTO0nzT48K5CAWT/gwky5BYKQka60xJqOFUynu3Pg1lP2ZU
KDCJg0QS6rbkD+Kym+yIH+4L5eMTHWZy3Y0Zv6kCL/+YF3WqPUXPPQhfEdu+LfjeOd7lJvWZXu+A
gOE9tI0jjOLJMdVpJwSOAuKZinkFdTNne8QICUqfwGoxXndPsj2ZsnBZ0deXq/tsMOIxZ/Q+Fx+v
j5cG2miDED3aFJkMnZP1Hh3bANWK3T8f9Qbpe+5zX9rHnj+SRlEtN/PVMA928kJYUl1SjWUTDogD
FjoL6xdP408ZdXUiDVCi35iPhoJx47rhx25bDK3fBj4OeGURxjF4OWmZckN3s7rf6tij9KzMvgEk
Lx3UTNTqT/qkFKhcMh0zuMYp+/Sw1NI2mNlM8D5KHY/wOWnUdK0qN97XaxaKx0teoT4usL4PaaDj
7ashPrIjaVw5AYq1R7y4q5Hm7htxIwsR2ms1DeC4nqf9D9MVsaSo6n8FOLZXulLTch3y6DxAhqG1
vBl4OAjMTtwTId95JJyEVZDZMz+zqsoUVuMpCrNHHv+XkEmwuiOwGNsUAFIVKKnFIN3DQLjHjelB
15Pflypep18exFqZBN3j5GPkzrQATKocO6KKL1bDKNcNpKiimX3FhRK8HLn2D7iY1vqrK1QWfTLY
4U+SF+x12CjarzJ11qHMSPFzbVxOfjYWSjV2F6oZWzTnTUtY+iOq8ATz0RgO2++xmsAdUVspJhfT
v0o65/26GlI4s/by1aL48572Cpf3vDnQb1Dws/XFCyG+Ja9/qzuFhEPfOxBiLSzOPh/RK4jcWMvF
9WHt9c1hRAcXBSQe7922Hp+zrKitdOLP4hIuh5Gu3zCs+6eoFUiIAEGFdpEWGRB5/jKZVpER9bXL
eXO+31pFK67wLJAmbugRSrqC2w+bUW6m2JPSUtlN9ZRatSe7pAz1xZHqH1XrAGGufTQaK9lJr0oM
fgqG4v8keX54+4ZkQtt9y8XZZzk0oTAyMAlytevU68xqSdwBeGBSVQrPyvoF0pItOt+8mrvczWL0
i1FXJ7mimHWbk5lXhTrHIyIjfr2gMyzvm91MyKizq0ZBgycJ8I6VoUKc9nC9R6w4Nv+SJOJ9DGSv
zAMI9rEpA56aJvqh4+QrTL1DJY/zGf/7Nn22QJysD3q+lT8hcjaZOTnzk0qUb8jzAiosk6HQ4Pc5
2TkSEmeOfa7c4L81pyTw5w12FqA4riGfIVr9w6u/LD77/j3xIdrDk93oX6Kh5QpMaEb6hDb5NojM
O+mvAM/0MPkIgmNsMJEEMuaZdFox8EuYEZh3xeK0duk3foIPKIqIDex+v9x8RfzyCa3EX77Hk+y8
zVl/wsZsByDp2k0Vuhy6tTUs7HKaB1D+S9VAolkSsQZ490fi3uirvWjjpHxu10ieYOjCeqDYyxwZ
9LTqTFt+t1+dGlzVPksNSCYaEgHbEqKJCIIXqHRZRL6LZ2ClQa2+npkseocn2ctKQbE1e3Z//QBD
ZyPjCfHdIXRlK+Xh1bYj5+ZTJR+TANJQWhbenVrc8GQjhwNmx5VPQlVkXAkjZIVYH0kHLhnAeiUU
LfAVv9uPHhf4jwIgQjHArp2Fuog5l10lhuNCkvwOQcJd44Z1xdfpMWKZVQZhl5tL4FC1RqcUr/0l
vGSPsHAkcDbiTuKb8taubMLeCQu4X+ByqW3eMpeBVbqVHgjHGQru5kJ36Jlw3YkthE3/6BrvxkNJ
+kK/eSQOJnp4Nb+c2ZFqxGR9FKkNmCwBqZdRAWhuE8Ipis9Dq4emwVQgaS8dGqBZ+Cjb9Hih+H4Z
KxsiTrullm64PZBoZpyib7eCfysup8ge5zcZqcCgCx2GrHVNM1b+glsOcOoerFa8bMBRdsCWI4SU
A7wFmxURYUaXEoKpYz2JOn1YlHA0NNfipFv+GxHMI1ovLEocohRHKm7le2G8OfWTkby84S7Nkt6w
mF/Sn1EIBY19YLL5U5ulzQJn9/bZxGUjDmVeZaWXe6DFx9imdgGXAJ7NLQ51vQqxUhWFHKsStt6k
Z6KGcGsRbjgLL5S+4YDV8UReqs3xaSbKnmgV20hd4WnGU9FZ3hSRjEnmIYjupgkTnDgdlsJ/8rEL
PD4lrPAn9JzB8sBufAO7fC2tUwJeJLzotg4AtEDYor+xU7zOCGSNzDFTN2mUqbjf4B2PAu2wnymB
RF/jOUGAfSufw4Sv9KByDhtTfGC1FldaL+S8odN3IH6IqKCSxbxupOqDRaxtLFe5Hh0ZbH4XGBQZ
anLI97LyIjkWJZhph1m1OFj1PIZOAJO++nQkNjv5A/BhxakZd1RYZ7SqY5x1obceiO6cbrQfpIHJ
jM6bymUmB86bZBfvLP0rs/p/eqKJKSyDhE8pEzV01/Efvr0hJ+dV80K9xpPBtkEXlqXovuLNXF4L
94WGnkVW231dTjNa11uTx3cQBB/uGIWf+N+KGnrpDYRjyHHoAYQAQrKRYWt1Rnx/42Y7Fk9k37yY
NG3ovMPze1FdnwsgEOYRWx+zbRPqCncIjoH2Kviaoin7D+xtc4R0oiC9DkGXrBdJIaYtQG/64gMK
zc6ADGKmPYq84DWsS14eT4vzg1XzdVmdHMs7VlyxifF5cfFenu/65g+Tn4DgSpNlU86LhVETebQb
4oM4j9G9Jvk0lbDs9hw+P2k/YTLefkNlEYMlJrw2Ie1IZgCe78BJugybQlTPRd25wDYnB4dKPEVI
ulxVfgb5p+kwuyXuxqliOavAcSuswUZHcrcg0VfXqmyQ9xPymDEGR1Ou4dD8rXCo+oPpLiZjhDqs
FET6iVbmgqah1xDlNQ72z45qQsKDeibYoZxxCdqRjLixSSg4umg5vKIO3BqJkRbXEZaAsaPXO+yr
xOxylDMg+jG3D9N9a33KFr1g7x/xpoXBUwh8O0PAH7LKPHDOJno/+P1LNMI9EWRkfftNq/jhpNhE
itp580t4cGPyPPh5TNVdrc4yIG2OXSIJLadPF8RnT35ymc26unChxMGVnHgCDJMAXEmrERa4o4Ch
aUxqCl71IQXEuLkjAdXeEBG3DAevRpUi0zUZvjV9iUcB9ilrjw1XIZwX2C6vY7/HoT+Xwws9Facj
H1EmfURro0xqqcHLgkeUJoDd04yO9mgprxitryVKqzVntT0HCeuGXkQk7DmvAwPfbANOrPf2/zr6
inOq4IQZPfC9BD10N5pAXHqBZgLHfvwVttzkVXUmepbK0ptDsvQy2u3zyyq85Bd3iKG3EBpUJj6q
vcSCCP/eVDpJTh1sqC4bzzvRrnsuIZyw330gEOT1fWbiZQ92o40rpnm3MRGQzk87Npe6JNQSz/cH
OkbawGXMDfMY1+eyA2UPf2yIFG/JGoxPoLlWJcOXAABj00T6ALw7IhIWpoKnplJJe+OyYK7qWMgA
WW1go4OQgH1yNNDWjS1fkneBUBjMFfBFRgTMxlxNQfyLzxIQrvFHB8rECuNhnndrOCCn1PHefoup
zGB5Gl99eAuvW8QDkya9TcSNRdDvHFKfgR3jU2TGLOUO0tSwpoXCLJg5pmCGjUUMDVqPWwBXh7e6
ztyAMyZ3OXI7plTrG9hJw70f2VTajk5jlRXVBeR8/V7kFs76EcVCKPYeLg+O7z+3BhvpLexxDsVY
RTPSNKt76RMn111NnNeyZ+uee+cxrOei00kbS+xU+elNJHoSGXVyK+JFkPo//uNNFzmnKO940C35
TowaFlGWQXhaSQOYlD6voKmBi53oBlOnSTZIAN8DUr49Hov7mZntso9mJT/St4XLeHs/w1O/81cO
gOQKKi0dvAJ/0sxBuajKTBXlEnyCqXDIdHvpyKfnf2mXc24JoKU9GFPI3FBsAaXfbMryN82gV4/R
Wo5v0CFv5ISxnBGADTlDm/gwMUIZn+50gar00nx9epFh1XX3LxY+5NZ2WHBK7Sx9YxhlWFMgOuCm
dhBhzQOwP1uCTknrAeiqRo1BRpFFht+RD9H0BjoHx9cfgZsv4GhxqvcEWJIXdXXq3uGIQvdPzs89
KRHrAl5KL5Dgo1KcjLCypBSl1kE1JUdtG9MWwEwO1V8oU/xlOIV/Fo9C/7SGhgnyCYKv1rtjFjYC
a61fv3/nDR5MpCNYbhRdIdO0CaP6ovSuMPzZkMdFrwmolck6gWV80kQ6ObRJiW59sN7v1oL0N8kD
8EGb2KcgV1CfOUJUAosZe6y87eC5BKRoKJAatWfcNFc8Aca8AB8SfdY76F1utor4h1JcKiTC4hqu
YTwIzvw7+GADh/NQhUHCgKAbLm//rb36Y1lHJIgWRYmBgQ/eVR5SzDF3zv4uAcB/yw2uI+6/Ht6f
RpMfxcf2kZdhb2yfnoxRFSa2ZudheV0t8GqRVSdws4FaiCiTvqyTy4H4wr9wQnLhQqog5EcTP+el
WaWnMteWKJ61U3iUSwcLV4JDntWqz2CKo1KGxkbpxCmUmXfDyi7c4b8PfayH5zs9VIRb5yqxRPk6
V+Nk+J6skZid+8QvvosQZw80MBW9qkcQMP3hvV1ly4jAq7KS6rrcduBcH1iS57UfTUA8DwAEWhjW
RfTLhQ1dt4glI1xxcdbKShzOAgvSlhONEkReEYn4H24lWsVd7M3PXcjzS/9d5FuCl/pf23sue4Rb
wI7tzj9D3BWDvLLcD1OX/u/+U6uDVDoGyYCc2cW/fdUZQ+pwe4shd4nKWLH8Pleh+d8JpYhZ6p6G
879dX7XonaDLfrAmPaWD/akIoQm+RxnE0b1PG1/luwYxRErjrq8nm1YYBhWkOxz+gIXuFRxDb8j7
skfVYflDFnYwCNh1hqJUB1DsMfeNtnxrUPzTcSF/FwnJuyZ/DrGBZbcqBtMqRj5m9a2D0bpOZcnq
s39SFOEAphPS0Qm3QWQBFmI9goQLlFH6kZ4UqCma8784kyDtsjZVITEEPpS5MQ6Z6+MgMork8Pjp
6sUEKY1L21Xn8ivxIYdenUxhUay0x1WiWmzTJ5kXx0gYQDbyRRSlaQhSluJG6TxmoXQvfnqGtyXk
38aD0feNQghsHz6UBEaqJwj8HEHeyTBs4Ou+lVM9WFpOTXaapsQYg15L3BG+LTObhhStNpBHGVTa
eHY+amo9Q4qJf9Y1HRvhLhdKRXJk8yXksBmuPwM4w+/DnfDufaGJmJ/ioYfzEOGPErPJN84BzBjH
zNbHyS8fStSPoPjAyfkY+U2FrjHk0+ueSBCBWlJh5mZZcTb0LKp1v79aUvKG1xvOXFY6CnX3p5YD
kqbK45Q3gl0cjCdKtj9PnDul9D0lgpIh2f/K43Qf71G2EQ6P1+Zq7HhSR+LmzDBY0yPu28xHPMYL
V9PU5brFYSiPJdu2MTL7/F7tyc0bViAwuplWjj0rn0yCvMyLgSXiufaGBxNcsVQi5MG7XYyWeySZ
4H0dkrkptkP0j8MUQG3EiKApons5fTAwrIVkWPZmElg5EQ6GtxddikgQHYTUK8WsRBHJIFkBWc1M
np5K6GduLjQAmifnGnxoisJuYT64gRvyXvRm3dlW3KJe7G4cvt/MN2TqJFLJzvEtJMoJj70wG3d7
YWwlTvqNz1JxlvxMWLDklHO/HBJBV7RcZoSzp9BSH88aeuzeQcjLS8Hvo+Y9qajGx499XNfGWJ1R
9eqX6KKhfeXhcdbnn86YLp/94OqYpAiBWJPaFa/acs663WhFL35ZNLkTO8nO3ouEi93C8cIXVJIu
WInKeg8NIW242ZQMwjBbtdPSKKzpzgNn4p+6dSFm5nalqeM2pR7X7zIjg+NgFtj/MxU/x/8JK8p1
fWxHRxt6zY58LJAjluBNleDDjOXEJjSAxQh/E+9Ds+SJj0Bh+7Bi035kQGz7l2NXfiy7rQACy3cZ
IXi93RG3OP/I9g6x4dXjKmdPopHgS9d/M/7r5CZdcajOKKQnDuqlD3p+WYMJ5nUszzqQMLUGZoG+
Fh50ndZt2eXrrDNkbV2Y8OTSXhpkb0p8NPOCAQ2VDvufpD7btFPIagShEo+Oshiem+B9nbKLbkFz
DssDCxws9K1p6EsF5S2yojEXC0fWk4IkEUMM6MCUXG6HP8pycVZXtK2VWHmznZ0mrL28k5aXiHyi
MCMAfmHDk26xvHH3/R6t/kqed5HgQd+lGyQ/XEDMRxGSxmav79jrIyOmo+El99FgpA0Khn8vwGeg
AjjEAKfvHqLNDdjRBBQhGlvjLqT84vRWmb0bMHi5yvqr5VW3meCelK1bdzzTPDaTcfWu0lChw/E6
h8G8LkcXLGsz4SFsF/FToALVWFNFuuqiq/7p9MLiG8JnWYR5CyDY43cYdqsR2s0dqcH9Kn0YMToX
NaCim3tTeDFE/70jy07O1KGrOMMxwdCZ2kw8NUFK9kjX+jsj53x1NL5EzwElGdUQAsFAewVQEkF9
dKtSWZIJkA5YnfkS5NKPpDKioCb9eu5g3UmbkmBHytt1FetM+yEWiA5QOuMr+QDATPmbihoYwfdS
R7qMdD3DPp8PbUC/IvTlrDTsYz0Scm5VrCEl/x9uAbidRscTlfMVjC5LWlZlRw+j8MN76gW3v3sI
lu5HNKo88kEQzLebHajytbCJepVdQKuue0BV3Vo1s44H8nNSCyUbyXojETzabVXLalipLmTxqzIE
ULSLPXfBXzW10yZH2U8IDQ0XQyrZBabbKGR55144pqeXK+eLngEiUvMkwDKHaCclGS7DJIG7cu9X
+BzLXsmXZYk81JznGPuIZREFE7NdbW88+46v5+tVDbrTvMRTRDqc4vnCMUL2I0Y1AuGZFkN6lSQB
IjuCOSFsYiJXBAevJwDi5aQ+kSmSgjJliXuNpcvMuXC6nayqxDJynKW+zXpsrdzIkfDex2LBoMxh
efoiDdhwyCf+Nv2IiU1DyznY7pLLUA99C7ckNOLmCMye8V0xwT08a4mMnL2gSwwMtL/DsxdP+Dqr
YWTI1W11xFH0DYPKDkzO6oJmGnouE/mWpFjz3qE09l9wcgI1x5Maor+iVQxpvM4qaZFNn+GR4nGY
7HTKCLY59IY4oujjItTCDRYvcwDmd0isdoNZy2/hwn/GcbGVAPOkLZlMcL+jcocGELPTLXgBI96M
BfiujDTTH6YxrlSz7H4E08/bM87rgq3KEkk0AEVC337XgZIgxmZpwwtiyG0xLhsSp4iaF1qiAkXk
YjKlwsBQe99yQOlUsnXgfqGM3A3k70XCuEISk4uX5NdAIiyo29u5wzJAriX3nXp/fThxwHbjtuaM
dwBQDBAcQccs/5UMXQr/0ZkTOwAiEBMPI1aJ4KDVmUcBYifp9YXok2phG+EjT9W21nmg3NQVJEr4
6dAvCzW9E9T2n8V1s1U8x+OHKTlWhqTXUA+T4rGrvNc6LXMZ7p6Jt1eL/zjypoQg6EtzuqZBt72W
SNMW1GGMOYn/xk0978HlRBGEzD3/L7R678BXGmxeRxtr4UdcAb6PXMK0lDpUrH1rc1rWXmVGS5H+
O3tiqkqmfYvcbkaYFkhRBuACpc6mC9ztHde4thhu5zd3TKTxKir8Oy/+JrzLHzC8Lfj1o9AhQ0VK
vz0QfPjyLwGUM16gRjVlmX5222vgQy0w66L0FwjxeEgTEyjjTW8FxmIPBp39PqyaeD8XPL6vMy8D
3vjJaxqmCcGwQDKV0JsoIQV/j/edDvkgeYdV3b1fo5+b/ouABV4mg0oztL0LcOyMWErmecM887jZ
uYSkJ8QHFw63M7S4kPTWLsoEoZzzMdjxTNK3/q7eblbWXXbvwhsvdfpHXnE1WulOWJnGUvG5k6hv
99ETOPsLQmPK4wZ34iW4Gtew6CZnCcwazVvuHgeZ+xPKGkZT0YKcDDslVVl8gAsK2hGVcj2BiCRI
ZQx9zMhfpabWqiOhcKogDgDvlAd53Xrs4ULZ667J5QGnJQYKQfR5oZ7jp07+vo5gh4qstWySYSX/
RwBH4vTHZ48WHbmQNV63iEU2AyXpV5fT4PWYeDS6BM3XOj8EdhSAfIw4KPGOY09UrS028TWEjyle
tKX1t9F7CyRIQCXlRaWUcQjkxayL+1R2VxMvYvuhkF26ZRnvBx3+UY7z0rAz2ZOe7wAEMF7b0Llc
rz/ROr65ZN5/IuDMj8ioCAFXix1JTebHUEEiFjUIUM5SnidyTOPUr+k7GOACGi44TW54WXVL9XSd
j4zPdOHkZlF79I5KMPZdKQWtJ736sLimZEPVC25VcQ/glxzcrq8ZX0SM32WW8bKFtvyScDrQb2Ti
llBWaOXDbSignJ0OFp1MXw0+t5+xf9g30nKZ1mM7QbIMx4q+l40MHj5vLdMQNp46a6diU6SjSFeR
gE2SQqAUesk/HLUJwOPkO74a5HiG/7wr9IoQwRaN3A4isMB6wFs7XjDc+yxqSGpudU1AYEZteY4I
MB0LDZGrOYeBzHU+DV0vG3d/Kbjz24OHQguLkru5drGZdNinSkOSxiCDyfFTybrhgSUpFTnhMCZP
hTzFvyPi7UXxQhIupDmGDDSP20DGYv525BbT8cC4ESBLtFaGa0m5m7PCUwF1ubV9gwKJgtrKSwcU
eq13HuGKbGsAHjZmr+Jm5JBRfWX+kUUguEKZVhF4I3cQBTKYij+oy37T+zI4+zikCoB/P2ujgGQA
9VEpR1ebl2XJ1d7EXlGQYzMxBb0rnDOHaOlCBR0ywA2EXlIZVEmsUIfh/qf4Ca80nphY3wERgYjG
1a2oHNXcRHndXm6batkdJUaWbr9pcnWk1QHw5eEqJfHyFeib+Cx9gJ0KKC5iItBZbTcVSZU/G934
Xl5AS8Y+sRr9Sn8qJxtuZZ95B+cszQKyxh+tsl3l4drJ6mH9gtZQmkdZFk92qtQTqRAsT6ff0N4B
5qmTRpQ4ZF8AIKKRysCPDkzRJcWqTgvYYD2p3YsE5iGVTKBrhu7dwsUhP68BMxkE1vmb9CK5lQck
ylGPU8+d9uV+yz0u4j5J2krTDz0oe2DbGVSMLAxdKInxBPaTLtxYY7V4rhjWtg49Fo3rd2d3o53X
sWlopUP3Krs6Z9ARaiWz/EmPq62hYB5H2DnVXhUyUjoqJPrMFIw1XjaIBbJvDDt8irHvsMyZTDXb
BbwPfacwTLrpsMYBgfQhtbuziE9bG7qjbGhZPLe6RugMAoFBMzw03EbjQoMJGiP9Ug02zA8l4CYS
bGIhnLLAIpsi0844y+dMwP+07zdzGEzJIcYklt5dxL2GllCxlfr6IJyuUyTmIbq7Hyu328LxDqNe
qqAvGJu2bH5tr9+NVxecqL9NIXn2PqAKcz2Aib5fuAMbsMz2TDb89OWlB0/iX5zwuegxEalNkvad
bO8omQ/Q/o+LY4tQVdJ1dBJ3k3kDya0dod8JDVuSQL719fzTrGJc5v/PklTkh4NNOzgUHZ4LLnM0
OONBdkuT6VYWG11Pds92PLtSMIuitH9SSqMSaTCaAQxnRW95Oae4JhOuWBayyT/HuyB338fjW8P0
HBPPCWgnX4Y+2RYxSazmLxsSbYK9vUzd5mewNPLnUyL30Ypyz91oPzu9XsKQp5yCG2ehHAROR2cv
kvIWG5jg2cRFJDJbH4puGckFWQ9pJutXupz7tnd+xhY3RFCXbRzMLqJovzj5OVrF55X3WlzsVl6K
QCiJfTiMCbluuOxwRdqhrGhn0qNucHaMhovQgtTNWI3cn3yAJOg00rEGA1yA2lykvadBKOpJwovM
ZaZAR+b6X7N4bbsvXcj861akY7LA28A7gXsFDVMUeWrJVHUvs3EW5Iz8GuDfG82TbKYeNbfvv+pP
PTv0Vz0kvjqSd6hi6yMNK/+zWaXq/5nQHfBJSYx1k9hL6RG/5WyFvNhUhL70mCDqOAMZmMafR4XU
QDUhxF1EReyMBdzQcOT8uu2o0zPyWx8Sqln1319wIBD35pw8qBjEwMSpA/VV3DLXaOq0+tFQOXhL
Lq8uR8xdANb1+/OAiITq0CiKfbBrZQyQkkPgHbcYVIahjlf9bHtJiJIMM79mla8CAnIKMT8QfxfH
Wi4XDUvTlTXbpfGcj5wTdJAA197k0UuyRvhBhBKJi0q4wTy8aTAAQj8kRCMdXe35SagmkwdJUOJl
o9sqF+/IyO6vul1jjRGHOB9EjTw4+pJ+kwy8V/oPMUaA7FrgMXvvsyzMtSzC08kQ3PsLMJ3z0m6v
XyqiA9giioLDP6HvtGI2TNDjqxrOKKzns3MIQGjLUv64DQvAzChcztT778aK1i7eecZbLDnr/olg
fJ1WjAfo+1Q2l7ulTNGBDG2r9Rt/2vjQ9XyjD2pnlm3ayettLBifDRCxQulhCSgiS4HStT627erQ
+KNTUE3/ptOU+Kb9I1XMwU6A10pFKE0uHVzALJ7NBO3BFB1OkR4Ugjxp8qdRiF3Zew3SzMgx1EZt
aornp49bahkEE8UoX2f5l1CXpDHvlYh63j0cC75qLpaz/jIZ08EG/PZOB+YyqMKb9puqDer21Tlk
zq8LuCHcSZhfduRzVLlf6+k7T4ZQiFUXgxV0PnrH7yPsSJMeWtqPFDIAXx8JGE4sK/Ja7Esbc01z
ftAaigIaF3f53MRyS7FCQEK6O3BZaoIGAc7Dklj0NIr7YaY6JWePZnMtVxQ+9apb/F4C8VaARR+4
J2840iDBj81pKminFjWxtdJ9nBseAqa53bz+TJwXiV2XjZovulcd+QYJfa88ROmu7mMBcqfp6VID
4cZR8jpPEJJcQqysO/iuWmcJDF0boWL7InhYV+V0dRo+lAWLXNgIqb/o+7edybkcLNswgHXNH+lz
C7fJjKcFak0Dr2+ldgaS9VNOp26f9V3FqjwTLlxIbZIKWLTJ3uL6I2pLdtZRLo4aiL7CksXGNpQ0
NtGukobuPCkNIbMUEU2Vwyjjr5q2rqkB+oDSzhhYCByHAk5EusXwbMxrgJICiWBxWF1Bu61XppLP
fdbstlJPn2UDrzYJi2ubUqVqXmsZRIBwNyv7psYiQMQscTG6nYXHaB2SLjN5MJczrIcLAjlUaA2X
VLpME1ScaENt2+IdEmR8a71PpYTXKUiN1Hmdwf2qEWx0u00AZe4umwJcCiG2Vp/rMtfOSwqaPXhX
nHGKBdlLONoIuEcrS40KT8QJcKVPfMy6uXX5C8XsMtXWbyiIODA5/BLpX5/UTcoeltty00Czf8pD
E42lNg4+7WPqq2ekp/OPd1SPonap25+LPL0ywMkx8+ZFp7eOUzetMQKtTYOnTpalIc29sHRF+1is
eVHu9ctm1WTTjsD8CpDjuaTcFIcfvWU6XkSWYVlGQmT6BJVexjR2gwI4XuNDcY4OZqvUjaR7aSgI
dOMOU9d2QCps1jK+HU2YawbKpzscLf9wjo3beiV5KwgvdgFK4EoxQRyFWuopndogWVlcsZkobJY8
Y9c0PE2MJ6lme+iClyaSGy0/Bu8Q35k3brCRQmxno7s7KdN5SnIKmqulMsOvAElN5qfKYweNYIEi
Wt1JNSFlCZ6xLbA3g9nN8sQIn4v62iizZ0NpgnhQHPELLk5Nqy8XVOPa4eIPzeJAJ4gHN+4jXkpw
EAsf7ph4Tr9rGZ7ZjsT9WGkTdYvKCOmozb+glbRAAGj/S6rl5dcYOh6nujDxdhdD+JbEV+OIum4g
eLLoS0HDwk4ralohawNa8MC+vW52WvmgIGMyfq5ehHCqUAIF4R3BWbEc3lvTz8MXtD/kpKgpUySK
Zc8/U67vbzHWyDMs44BXwpDIveGQpmdeFp0xtXtkhcPv5WQUuQxYHG7kdo1g0qOKgJuJkAZ3wPvA
UCJSgy4Heks5j8KHJ08OGiuX71NCvDqKIkSC7eWzVfewVpQnA7bVy8ZZCzFFdri/uBcqtHgrFwM5
GefbqKMjhLmchBqkxoDenBfR2oK+9PspBpyZLfWB7Mvep6gtfuGNLsSRltAurHrbgICC0n1ideIA
e88ZSkYNtcBIEHZ2yNYfgVOBaf7r0LzyvSx2q362vL3I0nwx5YkoQTho51jrg4Bau+jCmbVyTP6N
frFruXblNxpvM139iTb/aGJ5JxfoOzDWkidgnwl+PccdRAEtV1vAYkQhSE1WApgpyy3lHlGzS39o
BE9+9bBTnW0S7evRcoKUGYkgquyPEA465RRglE7cbJpyxq3cNF+7ETE2Dtdiq0ikmqpzkbGAqmd2
Lb+K8w95RpuhXMPy1w+ZNSXdDOc4WdRE+zlYgUGKtllY4HijwYRkZtIPt7H8Yg0MlGhQnTHNQ7oL
H64JYCNqDKPG2zAbsO0IE+h7N3J4ajPcsl3qD3t8ollvd+6oLAarUyjUKTRr+bGj7BMk00nVEX5e
95IUbPWgIzTbZiLX8+Os9ZFN0m1+jvYpZtZtzeOQA/PJSbmKtiKMQzuxcO3TNxZnpRz4dV3IpxTB
2pIJP26lde3qPwEmhMfn4RWq7bmegNHHW4E9gByqFYRGsb4cKQcvEqJWN3J96Qvm2gBHkwUWy33E
+eRzFbDbMWoYv/zSkAWwFurd+VWKzDvURTqOM9MGFtRGsNhAs6aaemMygb375t/ABJOyxEvH7eS9
KXLfe+mRF66wE/z3EPI3FztyZALtuAkf7RBCiOjg8EPle2OkWB0KDIFKZA1edaJ4IeWcLZ1B3YbH
vC6YrUbQ3aKq+NM3ny0ioZ8zQOUQrQegmvpLsLFH9PDCfvfzqBm6/FlMNKVxAIKDwiJLDx0HzK0k
bGIB01wIl9nSy7BWS3xxu2M3Si2XhlfOppOqTDW+XJPjoKQjsOBIpAc41q/0JZx1kL9rd/tvyIh6
on+A8la7fXs2vUYLRI+7g2q/76S1NpJnH/qwmvko5iYkoyipX5nIoYQS/ZtW2uhxl2ZOi9m7t6H4
OSjffJmquNN3JggLJTfpHenWZU/NeIseLcyGmLuaFDwDwdkkJXGUCHH1ctZtRizf4kSkzdXx4CKi
riTxEG2hpI1B1MccMrvcpyTYMsyK+/fXvoz7GSdyzY6U0Zi/kVALOExZapxOtE8cOOYOezvNoMXx
Td/MJpEAJ77jaExiH2DICBWMygac6o2aaBOEvkosO/gyV9/J9wk5cG5W6cQtgj09uZqa5cZ6vOfd
Rlj7cvnS2CLbXrHIKq81Q/L03omUxqWQuot7n5lUYmpNPKU0018eY68u7v3AGr72zee26OO3Mpkd
YQno1PA3LYM0G4NyAxLgpLFJ0/olHu3TIgyY14gAkt5B1AmQIbLCCTosXuacorvhSXekCwaFjr19
BFrdNpwPAq7S4i1cb+5/1SltPTF8jvt6UaGZvcjfAeHff9d7gsKfy9hIxpTMpR5QCrGutAhmyets
dIbCbsa+c4UegOChCU7wh1R1pp/FqNt+T4hkIgwVame+HoPb1r5chgZNITie6f2Uw0PPzO1I+qYt
oLRU8NhRxbaIQTJLVtVQgxq0K5DJXuGPWNBQzZd5qytWzceNGNnnl6elsteN0ocIwjoHUMW3CisU
9eJt/g23lo8NAZJQRu3FgmbrVU4cQEIsrx6pIadbOP54fw4Kf7V6V5fdiqH2strIqGGyS89WqTRo
EGN+B2J2YkvhBfUSc5jV5F85nf2/t6oH11cDQ/JPIWaDzifWDZ261Z5TnnNQMtT8atH37YGSzbVV
m2eGcAnUSepE38g6LJXxtVktJJU8mO5tXvDPcL+KwHzFBkQY/p5JCbiIOtKMeifPB1KdECNaPUrH
lt3adlf9T58eujIanvCHVPY6jkKDzLWox4iJtalwoE6Tj7IgPxhknmdoTwUFX6FIEgPvjFON91HP
upjXFchnVst4JEgABPw6XlvjgTx+ROGIT4ARzlVFfCUlfk71Tp6vyiYSbaNJdiwbv7WtsgC2J2dr
lmrfGS/LFrqgQLdyJshKuLuH0C2jhulrNBSksCGIN0hhYpcPZbbVLwZvYOUfbBO9nKbv75ou44tN
kVXzsC2r/0Yq3RT5HF1O8ITr+mALy/1zYOtLjnmBHqGounT+NN+tvRxnvYCQul/tFsKD0ux4cBZO
B4tL7p+WhA+2f11t874U6PQ9092K5VeLZkwUX6a3FGa7aWi5tTAwgIMWdK0z7kQd1B89rq8WXIM9
3DMicvvSOT3VdElJ7c0aKRyG/DHqbY6B5L2F6Ytw19xST1DaCibej297gFnbiNWSFaiebv9j83WE
ypj9lX9t1AZzIfOZwZE7l8LK7JUOCD5aNrU/54bWvjLKFZgGXEReyJCwHSqof4+kVEo6MiUKVzrP
LgtSXf8GWO8J023GyNYGnhy91er4Pvl6PPutDKM9Ye8Pfj3rIBVi68kE8xeLq6AxbNhnOekvqP8D
kEoz04gr3UOPMq0Nfx17Jhu2qxLY7ypz9no1m2pLdi1kcNp/MvSi0Fe4a0f5+QaMA/zy8a6s6ed6
BxgJY5VD01a8xrvOXCSCt8sEpQ8y58fJtQU1Zc5TkU8WFTSm8312FzRRvbBxx39SYac6EckALR+X
XvOnG26LO9OWAa8Vb2BEEu+u1RPye3kV1FJ25dtX8yzjyIJkyR14sY+gCO7awkm26hwujB0dL+Qt
rbmuGU+2xHrMpe3ajGAhrVa36v8YViKg4l02IE57OWF37ErVpbaH9CHSm0Mft30nn/DoQgpujYIQ
WhN++LDQoFSZMVgszaGoGRNgXD96qIdCa9twzQZ5wvhra+Mj4LofbkIGbsOOc/IvVQHmQb0+IyOa
i4w1S6L5FzHroSYPxy9PQX5tOGUgbUeY2htpgtyd2nh55O2Fo663z0oPUUe8eRSDwUD1Dw9UJn2M
nFxwRTxQqyMhdf0jpUs9KnRH5pySiMzsFTZTqnk1i58YVvJHj+XdMlD8RM9c5w6+QJ/7fyLwjEKW
bivKrCNSEil02ozF3SPPkHYeS2bqeeRSlgxDyonMk4sVqh7SpbGweMS7OqcbeZhyaEPRJ5Vbbwec
4gmt/BFk2qMGwx5bpUid1YA5Y7qx4fAPJjx8wUI1p2+TuK/a/OcUegJso1dcwn1JMwClyZ/4xLKX
KxBD5kA8ZjsQcnVo75Uk2UfsemYjAMU57AJ1V7YHSkxGMxo0V2eFbTw2HlNyKthKkNUhNP7t3c4i
Yx1z7qY+tL7SU5WCu/sacb+6rPIYUkQPlmGYVpyvNBmNopgOy93oh4Ej5fuqhqZfTt+Ze0KywLzm
jzXo9CG3Kbfw360D1Ifj/K9Tq27l7VBUQDk6XiwKvu0ogc7bt24AVAUwsahQ4tBaE2JYI5qUB4jH
nB9xthu40etlD7qktMnJ8s7lpbpuPBkPzjjCLt/V00JWGqCILBTaAU9E3ZeUCzgv81EYq9RMyyZX
r9twt2l5u6VUlLX0aq45Feyb/V3Qg3d3//PgKx9/ipUdyaXUd1WAB1Js4aL/+pURgajcrcg7IkKb
/6D2Y7UmdHZKQn+V8AFJ1LCa4KpuVLmB17yKOarrNlimTNGqpuILdllY1k6gBu+2xGq/V0pXQQv6
ZOMs9Ar+GQP6tiQq0sA/duKgeUgbbdRKCPp4YUgKsuM9s89IyyU1WgTKNF14doeza0UdDS/lcMSM
V8azs7U3RykFvQOEhoeoKeNMj/rBUCy4zcYmE5xtEPHXzxYZ0japDi3BelyBrkyrptZExyh8Eqvx
atU78o1XE2T/nQ3IcCBJML/fF1YxRn9w9qkoQHM6Eb+abV56qn1RSNlmaO1+5bXGVL1SFOuu/or+
HNdFkoZsulLvdgDYr5CKmjLHGpV4eAur7lwt8vzDL6NFhfNQnKjtF0BijO5H3CfY7vuWrgAKeMn7
4D1D9r6iQqZIS43hWetHPt2utGa93+otr0ZBUmUCUYU46o0+8BHaZBQesQmS6ayThMmXh/f1/SB9
IGK5w7QFm6Ktt6DdcHhL7U/WIG5iP1LDy4gx4LDwyDTPXAZvKLmrLOIGDzCuQk/NVJwUNajFFGtt
OeAeXMAi/CZh98u4FBT26O4jhN1FDAmxrMampxfZXdHdhnboldM3B0xzXxBU4KARXyHPhoz67EK4
5urdMULyAK7Mm8Dv6/I0ztmPHGsMXmUYPT/DLX5N1TP8U7nxm3VZVn4aTGkT1+zbKHvvjYYxEnXq
UrIMg9lEh5O5Bae1uMjK1ecrDIdXrNOw1stE0bYfK7Os6z1LUF58v2x0dkAyapWDwNUuINSKkxV9
hBXEUlmfFLMUJp3r8fYKwfiP33xJE5D7ySq231yXGkzvW+nwnvBo8XZrzx9t20xyEUbT2KKLiUG5
BDvWoYjyzj56y1ukxlECIxq2mKFAwZKx6fubpraYJCVV8RcRHTOCrmfNLOY8Md+19g9dCAacwqLa
P/tUesUFHm5rDqUXbLX1yjRbEN7AokYdMwAagyrRItBMDXJyc4KuQD5W+baaIKDCJjevqA5i2O5D
pJThr0emg/fbLFL/wl2DlSpPxn3UBeNgSLT5996NvH84HHnLg3ayLrHtI2pJwibLmODtUbkHsQKz
AKdXw/gbaH4StHQBZLHxvJIBkKNoJhsFX/P38as8NM8BaD8rgZClb8BoK4PlOPGGrj1px3wECChj
LhrOe875iVf/Kh9oVitIzFEos3tBlZQHGzmhUM9DxJ5tfp7Dgiv0VwOzxVwf2fyBxXrstmv0B2ha
tnDH1yhkntFoOUpwEi4sYLdhOk8SexRsGLQpwIQmr46y55B/BFtRUUMwjRoB1DoZHvOA1VaKQxm4
kBSCHMeMwXXRiLXLPE1GYrByGq0k2hmNDTXAqPf1y/ZH1StaYrLo9JCKTzB8WOf4znav5j/Gjj+2
dOjXrW2Q0fcikWc/Uqd+TxptnMcuPTnj1LKtg/W8i6QA5aQclvJus+A3GQdlDPWsGTAuEz44ICp8
EqQuqCRN1ZK/X3RzDYgiwTwA2QIjVAFfd63RNQ0XbjVoq4B4hovJT7gA7FdYQWdbe36Jx/v67pup
mzJY1yFO83UH/26pRKIgrCFBUdKHFTAeV5slMGssh+uMa2Qspb8pMejQ3HP+s03iO+Gp6VoZpIDf
C//eFWS/p4+2qJ6Q9wI5xujTJzZW5jqi+JAnGu3ZSiaqX5bx8feWDC/Nuo/2jTpyOekNde22GynT
mSP3tnuY84KYqBij+Cltz3Jwo1WE9dsEnRzoPbcx+4te6wA7GFjTLsDSKdfpF19T2z8dJEwz12dX
27EpetH6umLqjbkT9pnpNdM/yDeMaRcKp8+u/jnUw5mkVwksyULFTcoezgyGcckUafIERzNqw/HY
U5A5tYIvsfZzcd+AUUWVVLsZvFN7F3VXEr3WjeQyBQPBfUUXuVc7m3+tnbetjxfA1Ev9mFoBb/QH
le03Coat8cBtwLttpJ4qpd9r6bnSnqMSgGO3mHnMqd6GVbgKKrEbYuXAumiA+yw2hoX2TQdSWf6G
aOZha4qm+B86tPL396l/YK/sCisMROBh68Pa5BnDMgu3vygLmVknW0wE5ExpUtzkhCIybUsNmSlE
1xUoIQZ/3pn9GS0102F7lJzLs8I1S0u1gPxIiBmfmqpM4kGM8G5dN0h+Ro3UBXKiky7mlns+XuNe
Y/A8OfUbDMQs2c6GSWD3//oJAmBkxl5GNgV+iPFWwSqQhvfPJYXk805zxUhkmWqhC06UixcdpJkq
zzdBWOF/MVzd8r5eRMjaEbontU59bgBIkYNGqLkKelEBby043rHcUZDoth9hVkcfiq9GnhGeiaEf
Vprzw54kC0dKiOfzxtL9Ln9tkOBgG/TOMe7uJepeEpdq3pENfNkbbg4Z+btdYg/QF1I9itjf1O5A
K+mJd0SLocT+MfXyaGEiJDkG6YT0xWWad7b/bEl1tdN/lDV8/iJjsHVmaGiESK0yXsliFHU93SYK
etN4hlFTIzP5BtSUb+gTZFrMdu6s8MDQDkmw51BjfawF1sjnIX/sIJT4MZtnaxOnQuChnEaDWlDd
7Mlp5CKXCa91ct+3xI44Ct60idku8Y8V32zsSasqBSbJdmzy8uKPJXC9mzfYiYjWMsxF6C3VZMil
b8l+NitTpN6Q6UBgOY6ZXZgK0D1DXWCatIVHAyWorA7h/N/fQYDZAprzTceNs9gpXNvp33uPAuaF
ljSi4DbV6suetj5fye0Zyv4/zIWSoObKM0QQRWn786g9MJt5sk7cXt9euBy9FHOjRcMJ78p1/0PZ
qwiJXUwUiTyR2Z8+y+mHk8oPqd59LNQhJJVDIi9BQfXgbPC/UzdJ9EdBQ4v2zhN0vfRTIbKcsV/g
NN3xdhxbLT/Xastki3apOV9TTjNLPBC3AZNb54ubzvXSoM8nCe7Id6JbsoHrKCx/y21+hjHPD3Ee
290kzqEHmT2s0lBDHVF4cPkMb+HoHL9yl7VbSGG+U6l1scFDi4mJBCQyOJsqT3RjyKXzqV2xOTxU
08k7RpCi3ZUwkEo56rCk/QIjo30Y8+VmaoGx3SJ2h0nJs9iFHSiXVffL1cou9GyCrQ1rk/aBU76b
TYw5BbnRegOv1XfpPu5ASra4aAMuipB8zmhZefIiWYuU8zOXkf1vc1H5WBjgKEWGgg4CMSy6vAxI
qd5s44Wrtn5amrmSzdAs8om87kFBqjROvlTnJPcY8wtSNn70MHALjMQWt0L78xr8/mEvWJ/Ju/jm
cIbvFbKR4//BGl1MGEzksCenfJnyDHUITex+CfAh7ashP1rZvAtoOISO9a1Zf+g879VoRc15Usb7
8Og69BSEGv3JTql/wdP5i67v9zvDXu6MWbLKggFeZ8TEUeAIEnnQfkDLdVyRk5I2kFypAeqvOUjL
nC+njc0p0r9vj+fwF0SA2n3866DXuG54xIbwwQAJlVxU6qG4VZ6i0BjeY2yafy/S2SzBYeBpBgVe
qE4z7R+QLDF3e+f2WLT0n/HMD5QCKS6hYRUR0mcjcyU6WHvKGw5jepTC+k6QHOSpYeM2UTxVkj0Q
KjsvAoeW3frU+U/teMpjWffAIr8FUWnlsQdViLK4DE7+vG9/gvKQsQ8QUSxrhN3m3vEHFNTVi25r
ldmuBnk3QZBsiKlvRN/xYxrt9AKGe7ns5neufCID/6Z1bjZFswSPfJFPdK9tkk0c8hm6oD34SFay
KJSmzVAvQw3UkdQD6qfOzVSkmFRuR78etehluPbYI3nf2Ab4d+J+u4T1ntLuBeOZoaEE9dCE2BpR
HhmCk9pzolV1dn/jWMKgZyu8FSLuruXtgjSw2zxNLrheNNcddnDW/8y0hcXcIUR8PZnl9V0vGP+f
fUNt5Y22u5u2Bd+5F171cPdsaGHunLu1u87HjTUbcYYCMmisM7rhxHUP/8yqnljcm7a1NKMfnvE7
xeQK2HzducO6QywbEt/eIWlrieAkj9L2eAunnZ/gClwmMNKfbSzcvEabop/9sR5NI3dHjnGyBktO
z0C83IX/GhqM9OrVVgFLX71K5yyoZ9xQZVZusPW1j3Jl6aQE9TmQIA8uHtPamvyqeXpE9kJSaMCz
3L8jWZMNlLX3elAgygR83geuDYWQJg6KID1C+t0McaIb0yzKsljEO4vKjXfdHiMUBmy1MUyVhXsX
b2K/WstLX6dciAESUzmIM+VMSXZYN25WwcFEsv7X8hke4+w3ezW+h9EaTBGk53arAdI+hoju+rjB
NGk9JCiCoEY7/6S6Oinm4nEJl1Py+h2Qqj0CcdiHwc5LbH+M7mPhjua8+XwlUE+s6G7azaVRJTcT
Bck2nI9qTfh3SrHPZft795W7MY9mMVt3hes8bETFVAKVoBAGN/GCiPdRKd1ii1e3ZAjGNfSAW+lR
Cgqe9UEL9ArTW5l2iEqA9og4PNuGm5e97tE0n9R3licsWWCWrE7kUtBTc3RNO780C760jMh93Hj1
eNr9j3KnIc8yTzLTxEb85zXEz+O9cnjrqiDHoDo/6ff4I8Ve3I48j302/cPITbfF00sBxiFDD77L
93RxH6QV+WPcT4TAsNnoQJHwiva+AEq5lZsdH59tBev/2bNCkg9kJLeonY0MbAVKvtO/0m19GImF
6SQ9iPsMrEKIUH2KEy6qF0/FeBCcPzUvDO5JzoZWuJku0dYYT+QgV0alvyojFrUW+uZ114dqC0vi
aaAeelGzRj4QWXBEYOp+6wcKZwMsbneEaDSCj2+zcWYXZstSfnxn0aJR+qhu/KjSN3wHD+1bBp/n
R0I3tvbpj82qcZfvjC9v6lCnLA/3Ghwwnbgqmx/ZLjG0zZvOo+/V6G6lmPgSCSbVlgzHC5iJGL6y
yCSbdMKeVKyMdz+i6D8rjS1gf8ss2o+hqHNJY8QaOZKEgSuSUjYHO8A9uEUnFONCDTpy0Pq5Rh93
fAVoJYQ+/Hceu2tn5eAkaWUWV45LbUi/Db/EYTDZsgPd5N4E4eT/dfxxVHgy5iK51qoJQSxXgHU4
S9FmvPzQ9Vj0FlLKSTRIIpX/bbT5q1tmcfAqQ/J5M3LtcMqRBontclxPQFtfDrA0R5mTdGiNfhHv
zglH309sLBbwuiN4ihhl5vdsIKp+3otjToRTY4KQYUCrKTo3+I0j5hJvS7daN5JNhBXbpUS+ALT+
nTh2ieqVscLFk1rNQKuctC4sjl3hqSDtH1TmYCW8T/VsmAe3bgNH/cvfDmSGqqeY/Hag3R2lhEpF
lxBC+qtnCfng2HvEvL8w6jId1OK3vZzwVNROcoyH7Wo5PZelo5OY7L5WDHbJX4TBpTCmHkpbW+V6
9PriP9onXs920lxmVeM+tarLlvajxqNYrnZ7wvS9QCHWpbLpbcnKd1bj+TmhKKTWkk8HxJJbWN3P
HWhf7AxQC0hDVtwA6VH2YfmPczoInwlrLl96ikxYWKB1pg2LpPp9mLTpoN1xCeoI6kksSBJ46/Di
nkhR/TU1St5uiCY/fDK0cJz69Lke1QnlBvoDA4SfscX8hq4sjz8k/aUq5aYfpCgsxOecemXdiAwp
zkzY+K6zwL9Bb05jTwqfTiqbovcs7RwpVvzor/RrqoZTLQQql1QekCqrRs7z2aPTcEv1wN22KYMq
wMNzWAkP1+fsS270z2/yASpHOxmtVHbtxtq/5tAjkbq+7CzZ7FsdOz02YJBOsp6a0J92BwuaRP4Q
wC/FsBefLl4qH7n6+VDgPAAu8VJzsUo4pVBo/syIJFBr4Oxk0eXAPNAMzxrHSGHO7cZNmdJmEtun
39KgXFcqv/NjFkaTrPzNcwQ3+wE4j/V+0gpy0iNHmgisODQgYfEeoNloievLlo98SFZ4K3XQ38RJ
JQqtJCqObEg9Y/iQHmhuFSOuI50EDdUVzD8pMRz4knCNt6cJfvyPkKzHrk+6kLLROxIlqIGuB8R5
6/UvDhd8p834tk0D3YuuEYojQMBCl9Zc3WcJjcAzLx7RCpmD5WWSA4+m04KEjrOlw57gnxKX+4rq
dNyMcmOEE12eD1Z5vQvQa44106oDRP5ORP1LComje+oudA5g6B9TDbdEe0Slka2qjOsE/CAo/pEf
vdvXSbwAz1SKL5zGjYr9XMk42q19IYbpmWAq6yzQQ6Sjgu5szkckSJaPStu8TDJthdbfZZsOUY2W
FtFiP3pMziDyXr7kQJkbHM6b1kpCydW7k3vSIgO7Swi/RNfQPyIibA/0RrMFvglRDpGWLrUX5N3g
MLFhEb0yMhJW9ASLIs7WosuJAou3liUpatLJecC9+FRrtWpsFZslD5TmOPuM9BwSKtnQpYjQRfY7
sYld1lotgVebelNic1zgvuPYh7N14gNsTyYwo98fMpq3OpZ9CS/yL+nS2x+ZldIuFOo98as5fYjL
uc1mbXI/6kYC0ljgdjPSypSxnjrE69DAsnBWZeF2WHi0JHJknv2V4IE9PQHa2Yuou1gcrvwLy9by
fBIsvTzEQ4HFR5B3R1CJ/lAqTiB/0RW0rGBfp7jWAS0MzZwg7M4xIhqV//BMska26aA8+0ty6Sdv
G+k6JP5bxVYExaz8QSwwpI+im4aSAhHp2NLX1BQiWobCKSQqxFgsm7hBBp0bng4+oT7TAIIWKoCa
m//eCQyvD8Fq7BcXz7AFB/lcy/Kj1V2n9U4vmOyNmZEAvjO50vpdztkrScO1mgEf76n9sNXZJ5iW
HOabdYsYCDWSnT+jhUQwgr3upt87BuT7Z+moWkOU1WGGFI4zKcnN5wNs0WBYCW5Zc/2vZQjuXL7F
IG2B9sIEaBqlj7nYcMAutN9jVtmngdCJ/DEcoPkZ4W1O5++EDSTl5IahxOmguBQhCSjWhad1zmNe
Q204J+we4/5HhnJb8o0nURCvWk2Og5K51AhAN+vkBXFPTvcZC3BuND+b1RFjCA2MK1nTH5pa91dE
VUDYB6uX/J/eeNovvO5cB9Tagwmz2TWIcQcITFQy3lrjjwtutph2z022u7uLK9w8dXOUOtVodZSB
foLcXIxhOkOcIIKLfyj7oqaaRzytKLSqBpaj+rGWBQ64cQb4aAisbvjkwjXQLV1nN/EYf4jEPLvw
2Ym+wIv5TqBAkOhGp5yYzwtxwwpP6CPBE4ofNq/AwnGAljl0UAdFKA5UMQcZiXP5SJxAudjzw/n5
EH0D6VNnqfrs3le3egyCV7mmJx05mJIJJ2/hOt0ATZvf0PTxVBUoCr5JXHWq40KZNi9JaYxcP4iq
jN/9Th0rJMB8rpa6FFwjTK2HB8hTeC070uRIL5kv07+Ues71JbyvBT5O/GAa9bz1f/B3ElmOsjxb
rbi8QddSM58yzPiKgUBBoBDjwWeyuZiG080QYqqiCMh2EcyF5skx6Bo44NZgm0cOEoGrDhECje9+
4A+bH56iKIh9ePTvQ2o9F9mqDj20wp+jdiJ9fvknGnSiwQW82qEajspeSqNR39ubty0pEZsuBkQP
ztgHWlLO7vMkwQTLzgJrn7e1TgsMyEx9PyODUeL/KE701bajjJZVQuCp5gRuAQa2DCjiTrFQnHLI
IiFpD5VpkhYHpMyNwaKNIOPHK1if4fQmRikfLey70ZBJhHeY+7Rlj2zzgoauLJDnTEmFvp5FGrxR
etVDV/2Yb/uO/lAKuKhAEKqf+e17zTdCwoG+thHAHhM4aWBBd8VuFrUQQipxc8a0ngBCzXALq0My
rntCoqCk97+Lzld0lTSYvuUTIQsUIhlmUBUy7V67pLE06enKDSWq4kOoGlwcxoQeK3PRqVbaqdNl
q+JIKAXOBPLzGBbaHBa8rFfSMNWBQr2pnj9ohDrG+IvWDvUw7GsyWy6GK6zNl0f8hu5OQzeGS/2r
78dhfAHPNXz+Fw1PUHGB4sDnL2JsiKKS0FqZgm0QMnLu3Zd+FnWWkPKiVB0Ji/DOH0+7AZeM6w5S
ZNe+mRqkeNHTXkYMTh0KxNc7mWoq37qtvK+gUIQv175h/D+n4L7zoneQ61PAatpyY83pfvIcb2xm
VvNhW3IR2d8tg/nkVLk8bRSu59XAtBOrtClA+uzXXPtyw/DP1syHYZsnMEYhKKkVemdImc8ayH5R
g0xyQRgW4b5mk7Kbdo/B5giTTlx285nPeqjxZly5eT0YmIYpD/Dq7gry5HiF5Ox2OE5ujovSPQME
+2uF/w5JRa//A7GHis9sCBhBpXywDTHesk11nJeSZXGXDXXddh3UUuIsxCJW5XH7r85Pldx5EK1B
NO8LGraANJ0wvF37qZhEmPVa5y4y+MwcVYkSxZCrHkpGaKe+OHbDZkABYlmE6SILSVOs5Q4yvPlV
FlZcls4+wl1TUfy1laIXJn7umRRL4PehwmS8uoNmxlbT5TjRhmERVUY32wjLyOSvis27jFF/iGnb
hFgY0cZLmOvuRaI/zTIeFmr8yd6aqiHGgKCfyFnRf306trSEBMquFLJsJqPTzAC/vF44BdJx2jH2
3oB392LpTscOV+TtpgQ4Yy6R+vBJ4u8n6bLnmssVl5LktZCABj317QGbYqnJN/fTfqekbnQt8fA3
EvOsRX7wkQT/a9vKgr3ycaPbeeg2PIFPQ1vXURRQElvr02I7ClKfu3gI0DX1YYGHwS8OpUN6uVX/
d5PrUXWl0Wus1zBOoBcrsNFzN5+scQuK80NRVyTRa60lv1R7dwFj70j3+MBhoHsqzBgAK4YhowbF
aUgyhlyBGnQSPhUd5jbGEM/itHIiK/DkWX8psYwS/+MvZjHOeovPKEvWMn4mw1GNniuOgBhQKJYs
qKDYAWioqMwMzmYYveAs3UVad4zhLenzex6/rM3c9gGq+OWbljlKikJ7Ebm+NcyTSK4cvwKW92RH
3TaOfOYyB49sqTx+8TPz+bqYwVVWOX0WyT3mlD3Z8TKU/IYcUymYunsUOXt1kI3wJIWmvaRG4Y3C
Ly5Lb0jx3sneb4gagjlV1ehDsU5nVC6vYm8ua56jl+1he1+aBXY/dK/EOvA9Tg8ETkm+2VhUjCJU
nWeBRt75enyVwPMmxn76/gkEO9t0MQ9kLUzN+nyn9ienvbSe4b8q2O/Bddgcnx3FdWWhCB0u9DrK
sw9i0KdgEszhc83u/IzJt3bwP+RnZROUJeha2ed1poeSWas43aftEUG+YC24w6w/Tz7z5qeH/drT
rXdwuecTiDzlKr1LuF04NhrGNvNrSNsHFYAomYSSWKlQcvZQn0rxMBAL9yyi8WGsxR+S73fWvrM/
xTNykjMyJU4p1XDaKBd2rhJt5SdWStxoj19TD76kVelfjADElKM95G9Q4b1+AhgFWW2IMtf3A2rh
ncLen7x31p6G0H/w0RCxyHSBmxb6nInu5OkdapHF+4YNzIU20mUL2tYkTr7kJwvcfTlf7dETxqFe
crWYYbR+OtjKrJsHv7Nk019Luz389uMlpL50vSb+sJuhaUw6RFB+ixGfYGcgxBn/qAfxeCU6C05x
/gDulLSi8ecZprHou1UMVH/mexfyEZiIgMTevNod7rqiv1roj0wto4pGE5ubUBy85i54gpPTQ9FB
G/R0srfe0UhS4bjyQ2awx/RnrQQR1yYUyvDdiVlaxIE6zhIMlj9NG1whF2TIoA9gbjUc/9wJM4Af
IUY7XGMm3eN1/ZqPglrfT9M5GeDsNKYZuWaV7DxD825PTgH22XA5Vhs0arVkjPPEddtk7Lonw+lJ
zOf/vPXnyIUEKVn0cmDLPdI2AoeikniGxob3J0pquZKCUdiHI9s6qfiZnNZElI7xoa/fn1ZVoX35
buCY50IgXGzBEAhNdAeKS8yDfcKgENNsHkK8LvPs00kqzImLOUUAoQixRF10BsR7IJtWWRKeiKik
eQOSeHquU5BeT70gDUf4pgp2b9R87aEh+LKoFqQKCHQDAh1CJmLbKbbUJb21KmycARRe5D/rXckn
0AATL9YvLIwNMXZcROqXvRa0/5Fke3bYPqXJvs4bQCvM2auLTza82YeBlcwBGL9ai43rKpbwcTkn
bNY5+1RFL43ImXtXlE0ED69vzvuFz9BYS1yk2n7O9S9jRn8QcRpFbzEiCAnrfXXySJfg1qEiTxNS
jk5yHQqe9gTIS6nU8aECd7LstBTd71jst2qxr39DXWig3n31LlEGV3Syj1cP0BxQvu3YERmD5kiI
1qyv/s323Xst0HNMjGE7kHgg3nQr/E9qeT67m4CeKb5EjMfqVZwoFrylCDWY/dp8Hu4A/cZ0xM2g
kB+0O1b74CpbLaJ7tfBpjE8cvaGsnQLkdDsQ8NevHDGAL+oDiKwyomsOZWQ/H513DOXYyPjkjIKp
ygb8ZiJDl7C0avzP5Ky05AKhBI+E17lg94jeZeA+UFLxNlzwbH0ke00Xu5dVB8S1TF+6MGqc0tYF
1EHNHeTUqkpYJcvyNkESyjbssB0b72ij2kfQMFcI9eUvwaTT4aDJkaIsLZ7diW8FmG5v+MYXq+rk
3Xp4kzaiJMFMZoeYR7G5WpUIISFI/K8854T3RfTT51K3ij8YKhnFCCaTUqScIwex9a+UY3/E4teZ
GW+KPa2k7KEsHvw4mzld4IKAB4C8iBCL8f4TV/Hov8nrJD+ALUSa1Fi1vSHlqySrX46p3s7cjSGp
WPrLNP49X6AKz3UloR5SUJ6MjxMWXqKdePU8BYAkyqlHSDU72b6rmAvR/woQOiVWWr6MzD7ZHPC9
LoYsrB0I8ndMuo+1P6UWPlTdwJk3O+Ryx5JMXsPS4XzcwPTfHCQIiOfgPz8kOXMNEWn2RoC8rYzW
/Yh3qUNl7+STXWlccW1w7yYdbe2dmCsU47XvKxiN937O3g3ja/DuMW/qLrd5Ua81Y7dQquAxmRTy
YTJdANik5odA6JVkWm4lNnr+Q/vPvcxt0xImDrOayHREESmLOCBONnMjFMIM6zSZYYvERwpyftpd
4Ge/cFx7c5UbIXPcsq8d91//hBZ3oDHmG19SfPCvcopFUARHrBBB6UBkNY8tzoQ+dvbdP7mwutOt
UUEDjvmtgotlH7xI1JKOz5P29OScVcgzOlTwICAlK9AHGtRe/SpRQjZKCkevVlRtPpEu8pM8B4ri
hsF5BdQct/fD/2uCSVAtSv4Ja8IRc2aIUA0QrC2SE6PAMN2VB8540a8tjWYGS8Zf7JfGPdIOC3wb
/evbixsHESlhUaAGvrOD8+9qnP+1GxjNut8SARITP7to/m+W0C2Gm9XUPK/O/dw6g5ZLv1d8/fYd
RZHF8d3Ie+4tclXj/1NcuUgDkfvWal8GghiGTfXg/E/fs/XPr4Uwj7K+2E8Pm+8K7ZJpTLIp8HS8
cvC5/mln4LtgRSLVClnd0JfjEZONCVKIFf9o2gFvuJ6r7XlGgq1Rdesiyio249mTeQ92ExAlDeWM
rRhRAj3v21dzA9Ey9mmyDMX8LXo2etOyGyhhRUYY8zn+ALJlwpuUH0gaPnwuP5nhN8zfJ+ZN2XEI
LCOEiBFCnFQZT9EqDhh+fZpI2xieDweD6MmOkY6vqt62fRjEaifPG28yZuviWGGGtGzmc/2AUKSp
AcaJrbj/keJF21CRo6bJAsEc4D7uAJhjETcmSTRLnJ1I0QPS00d7NU20p4CFEV5DAgz3R0xQDfD9
zBSLQTBpvID5iWfoL/NJdGbjrwzyl/i05VGh6QOiu9dqfR13z2yxATlJzkqtwietDXx4b8oUqDB3
C2D/TqMP3OSF64U/sFv/Znq15ykeCpe9YupHlfptzmXqBR78ViQps9oMMBSkH6I0Bc4SDoJ1dc/f
OkgnhZVD+30sdl2Vwg+aCsc7gLx70Xl0f2awqhDY38LF3frf+H2r84q+a8BrqvNWpEaDVfLNGPVy
r353o9/PvP0RKs4xHXvES33sF9bWyF6PtevBV9XxXcNYLFjroPuBhgIJrZsv85zwcLnZwgIjzri7
wXLb+4jR0sIeVS12t0hC/U1RUgsKHTmXIhN6i/JH9m8Ptc6ihp3rPznpBmBMPsdB3gK4sIB8fqFZ
aGFm7pHHawFS1ohdePiOwdzHxlcQLpnp5akMtAY513nm80dJzFxnXQ2NW3Y+IrXf9QLODWAF3YYO
e6FWmGzezKKMyb01Ewp2bVucBEkesQGk7PNWw8wdDgKS9TMwK7aiqstfqpk/rQ99nRQf82YfY9Mh
7BPPmZRqQq+7/nkEWhOQv0AmD6MXk+ruL/++fIpSzYfBlie2xTeL+2+uU/gf49LXXe7rAJQVVxE7
LsnVURQHlbI4laSKPwgfeXFooDOp/IEHPEby5UXYQrBNEwbE7Tm4PPjmr3/S8YO5xTGkk12TlTt4
tcr41EII/nm7F+kPwUgx7Ul8RmvS9iyf9AuCmzNk4/FGN2TTK9ciJjoo/yf+fUsQvqetzSXEVXcF
TVW1r1AK9uKLK3BFhL57BQYSwnIc326/abRR9fewC79/3x4GnplYKgN6/mNRGbDdfIJfAx11S7yW
hujsqsmGOKYTpez4cFoSXVow3BfUf7vmkcyYZt2G/Abyvyn7qUe2C/9OW/kf+78ADPKQI/E9diEK
dDGoRtHcULZgkfz5+tHuhwJsVi50mpuKGYO6waDQfp1EjMw8TmGR1NitlDCWfTsmJ7BIEBMJrQx+
2Y0fQf3usdOWIdx27yTYwME7fNUkA286nrpTYWV/3K0lE9xsaCfs5Las2BTppeFHclCsbNPTk6Lz
7q/6fHnK6HFAlSHQ9ShSi8fU/Mk9KEOc2CUGvGYnnSBAHoT/SzO/XxF71zERjhGkA3rLWGa8M+CZ
wYb+gp3YEzq7czGtEbDBWwXm2Ao0Q8a8g4BdA7JqcSdpgescboMASv4SZ/spcGhKPCA1yptg+5Ap
TGv4qBidnyLhELhCRm2usRr+Qab8CiyFSRCTqqMQsF8FuMR8gtZML5h5+eyhvLxw1KPAZhBRV8jq
A7ckF4X92MKlzATsPUX8XtWC+ak81DKsvQDq800V0i74J6S1Bt2N4NEAWQr21cHPX/His1G1TlSB
lMZYJX0Q0NWLVbOWrk5tzPMMxLNxvtLYsq1IjSTwsAIxXtcXQK/z1u6cKpxcGE3vRFlYvuQaAhFb
lWjeIOnW0gwhI+qOQhUkhpkx2XXAMzYimqNxId758wu6dVFgNAPqh1DtqKUYvS7HHHc/0uPQj62+
rWghbk4BTBQZeyYKFn7G3B/Z2p4FjUdswgYtWy0KCq42xIL8XbiyQTvBEGDX+NiqtimAhr99Yo/A
zAP+NqdZP7ef3OMWJ7AC/kJDJuyMcBOmh92ug7gGDx1D5pBuPjXJGTcBZ8FxJFV3cd6JwCt+WLfX
OpuySDyG6Z9CVI4AEJX0bY9yhUFt4RX4upM+5R8YH+4fM+PuAyqOKp0PlM+ziyxmQ68yIGP7FK+K
4p1mBoxyZtGDq/7TXIby+bwKeoLl2agx6Pt5SqYKvaDc1Xxymfi91Si5nrk2DN9mQ1M8NMGRVlbe
lMEtM9JQ9fAqedWlCCc9T2npD7qNdxuOza5YNgpbmzQpSqk/E1Axv0oe6KZJCirBjJ6Nx0P3k9C0
GdQtWpyHrArtQfxgd4EXV9gSobQ8QCWFgQ7w3pifHlvyNp/xAdjshHeQYG0b2x8rEAEBqH9O4OoQ
6ERpqpbfu0eGm1VXYpv+iVF8M5l6rQU+FhgN4RIB2uWKjbnovt1WeFt8cDP/82HnXwOsr7+x+SnM
thbCSICnK1F3BVDDAzOOWVo1ueCsH4wTbzOuCQ45vWH9LRn77KDFxhBGk2xkEQd1lsIK9xkxADJQ
QfIbp77pj6sN/3lBXvtY0IWsz87gJFRH49La5hdMY7ZrC8ce4/CHx9xeb2UNWcuZRYsqqgoFlG+R
h8Nq0NrWSbk4DUZSHY3jOaP9jrrV0YAS5zc1fuJ4FDtNHf36t73tagexQzFGukrc6G9KOsg0nHfQ
AV6TMWAuA3/2V7ZGdbwb5m1/6NMRMH7K8WQV0bC+09DfDoZyPkt9fcxd1f9fxm6/so6QbYGqA05a
p7GJ/MtHQG6vb/anS/R56bTibod82F2AzOB7MMKWVLOihNkclzdYLSx7UgoLmmWMmCpk2MFjA1JO
Ik2FZng3deGIGQQEy+yoX49PcjsOOS0+zBVdaABFy5Zh+N/AtvFrfQuftB7zNdWsEDuZkG5d2MBU
bnKHrT4+xP8veBdG73zFs2caQ5s+x2utXr+9jQgfHUI1aTshfIoCHb6yGEgkG+uZ4IAWjDIvrRch
93oa2kQ6hFySOrbuT1gynm4a7GkCiA75QfI9uKlWhm4+TMOAOh/UcEHYbi/0ywtmyfp7adclVXQX
UN99RlKLgp/L7zuav2N01UvQn66mraiT8lzpNxwSUQZTM1vRPny7qLfjuGqFRD2EBeApBQTf4ual
GO1CsXOX6XiEmFzcA+yqK2mXm2PYY7Z0rNGZMNv/5eJD8TPFqgw8lAGMa5InDeODGF5cSTl1pA28
6CNDF0s6EXaZNKJTsYzSu9agBuCXNhSCSZqHewGtYN7cbZAgb8WeL8iYgF/jxXKIBdUxx4j0AAmz
nqzo0xh/dLa1BWK+OearkiM0yU1P4oue7/fyG7lYrvgAAbYQzeNyfNqb9wGoqQmc9OAC89JSXA53
R39+uruHxUQ+GDhsTdiIk1tA5lGKVzwzz4acmxEQQxQw7xrJDckPyko9GM75mdFW9g7Wl9phJt4k
tJf6YBhv15vrhE3crFUVumj1uPlA/iTjVtx4tSjdVxbPSQkcnKlSIFSOuVpoCqK3Gzsn1ioEh4Wx
oCxPSGtaqN+G079tL44RrnhbHX7WFSLzBS43I/kq5xk50eEmZ8c2mxNcW/AESLNNk68rv6JEf3gk
HuAchM/2T97b+gsInvePgoRB0H1paiRbuGPv/G/5AqAGd/SvHRSrGft3l0RhhoHg07OrJpi8KFaf
MRB6XYJhKEHkHsfgDAhj3Bk3a2koX2s6Z8Qc5+1ii3exmUkkSuNb+QzhOcZSiEE+qwPkXQcQpV7Q
upATZxT2qQyJZ3GtjpIP4dE1DLilZ5koDOzrQ08+wBEJddZfkPqfHOFoCPqXSBuZls2SIqlHLHpe
s3VGywUMTIuW3nqc4rwJD3ka+muDQx3jRLM0dkyRQ2cp8Mw1VCMx6aoNJzcLOe4GNFSDBXn22s3m
Vz189OeeiQjUE+E5Yq8kIYK2RP8cTdIZwXySlAUN/Lkl9MlQcrzXOnIfwf6a7nxD0ImadQyUoM6W
AAmXRAwEcgokH7mqXAoMLsLLaGb154JkoKIXJsZvMTN+APsVtPux6OciwrCCYx8egbnZW7POhsMB
3M8FjZ+NH3l9HjX+HYnlH82lny+uwerN5sb13N0gEEWU7aW/wQI0N5nvvJzq1tDgeAnktDxzPWkl
DxBpnHGBPjJJrg3cZ3d5QxEPdIK9dUPoo1cqrW4QOwOD3DiVyqJF08NREa+fSslT705GCUCLV6LH
ypijNHR7cHgUAatTNdUDPZrwIesZ/DYbVRgkL1GAgH+nnUik9L3pjeWfA/+yXOXkH2cm7qsE35NJ
PPBJgjNF21azBIpucpub9feShJSqu4jWmDv6HwK0PY8w8Tj4tZTuqc/MSy0/9C32XIpEjMjfsY7G
GdEL1+rLvRpmK4HWTouJRrh/RnRN9C58ZQ0vOMFc6qMABbj/pFai3vG6z/GxRssI5pLZnhYIZy9n
WuC8bHvuLDOy/TFNZhqs0FHeJrzTvlFzTarq4VFx3tQAkNI3n/kdx1JaSf31i8Dl0fFJUiI+SPL3
+9/QmuqcYnFqOdumSN6ZDINu7aTQi9UsitqxSOFyVc8DawqPYSw4IRifNRNvcLL7jlmX/JM1PH4I
kt9ONh+0w5tOcmlsIDRNcyZFssl3oKlxLGShCdQeRV+x4FNJPYexyNy7e4XwiiWJOBwmc21metdW
KV6JhAYxWbmgskyMHnAIsBJDZUBwZC5s48JqFc3mYP2/9rjts8NOxeU2utclpH7grjnv4Fx8aC7Y
tiFNGbcMfp99LuAbw4Ig4WKTOtxUAL+XaZ11q8eYNuvQiYcX7sIXAU2GXricn0sXnj08feUgdTQM
V1Ro62r6rtKQ2J7JuMSZLpSFkaJLE+eIqB0B4+xFS6CAFgYgMV3gmcB6lowuic4wXhYSiUm8yrAi
jew4ikrFqqCMOzagf06ZmsM81M2lVeuDbd+2qESKbxdoHwDGqGsd5OHjACNIJovhnHhQpzZEUSUW
ZJ5udye7ABDO0lPfOJPJyu3oxTJ9X723X6jA4maS+NKF0wQVcwjDjB2r/U0LASRb0Z7NwsuCA+XD
P9u2naR7eJJb8AAs6b1965CsZGRhnoSAq6Y6FCqp6UNvsgpMxbSA95EnYMJSKGcLGNXP38sY4j9R
3+/udD78B6Dqwc1S8Tsesqv/wUzJFuz98qyFB9tqP0dpAWmFY/zlmkvG57PskqMJeNFSOsqq3ZC9
H/Y3jAXsEwnFriTBoc95jmaiQGlmKgJNT8M5K7WIeiXmksepsHk9bnNW7oIvyoenqJfmcKuT62jp
bwPB1NIMNtJ73cyLGWvqlOUGWv6myjAHXdrhH/6oR0/RPXn5nA/6Uac5b/NrDEqallHoncFwOghQ
jLRTJ70ntzfl3xgPxVdoYI47XUI73R26fIGOGs4wu2f9PKGe6jAxQKIWJo5AvK/uhAgupN6mt1vU
Kq1pbtUVyy1TyROXw0dxMFBisgj5GbGnprzyG01zjJmQGCzclOBiV26z3RWgEbzncIWn1YDee3dW
oMSg7dXGX/pJEDrkSZw6ZtIYQvO1J5GEWCwhwfQZ3+rcQcSJlLPdZa/6B+eNV2MfKJcCFjD3bf2I
bAZJMZlxVmZezRGHB1kWeRvrxKKIhhGu6OftU59wqRXYHzcz2PT1E1aLW4MSSLmlZbqawowDZRRM
uuNG/2gFLkSeWcM4kHFWxb4Vrnw2XnvCPKdIeKwD0RRSpzPV7gcMyT/FQr2PJqYjRKVkW9eM90WH
Fle53V5ua07IYwfVZRXsIE87ZWwYzarNB1abLBMJ1cfmwCryEo/F5ZotsePTyDqXJFT2be/qEenO
b6umAZ85Rz/ZxtOZiNecNV6b4i1ZceIVacaSCwTrXnBA98PpqUwkHfYQmhL03td3qJXhiGkQFIuA
iiJ7HzTsxVIDL71YYeCECEZYTC46Jv2DXKTx5HbPGpcLsB8vJ8EDfA6HkP6pNIZLZLXcRm8TyJTJ
lTRvKx1VfCXuaEO6+p5OC6s9anrlbTdXKd6m2wXcLehoh+c/5YHTXhjjiAoBU9rabp/Q/iGpAMiK
FY5JB2LU22QDilBHj/uIOCC5OJfX+cUS7yr4NfsqSs8s2Mp0CfY38aoOfGmaMapJSMRsZOGfjh2U
D2g68cni/zowysvr9xAilbzah6tFd4j9pmUt1fvUioGH2Rp5LRlXK7iBHQcUXoSl0svOWPWEq9DD
Nt1HbpysVZSp0A3D9kYVk6Yl8abxCQpIB5zTVq3ElwwGH879TM4aVv7zFU/0OrxGZFqFcM8Voj9S
Ca3uoxOSSic9S4WG/achk/XdjcCMsu/R5+9kjpSSaSAwMtILOUSkCwE4eNH3G3kvqdaCd2fYXMwR
qKEjyRzd21yVHZEvEC6YsSCngC4fn0Sf9rTtWeKkOd/x+5/mePeEZQQkcZlEwuxxUw4Mgjx1W0LJ
qYC4ZCO90emnEiaKJFqBR9bgs58NQfWITtWZSijclwo/ucRnHtnuVjyt4Qk4CmV4xG67qJygPoYQ
8NXAjDrR+H/50CvrJlzXkmmCGGe3rqH4tuAZAxZHSx4+DR7/jfMRcP3kqSWf9aSmaByjRdyoOUVX
AOLzwVEziACVAdl9suTVOtno1XGq0pi5+Acs42jFc/nD8ZYnWEDYCe6KWqbcR05Q+hHUxyrwUPfP
DhBLB9MEbdcchqtSqzPbWUix6DWmXr+rcicZfoWkBd8PWSoR3OfCgOMbk5PHG8R+4/ivEjmYKVSw
7RNVHnaNIaG5QYhEeOb6G1kiaaMzfVVwKHGcTBlmcBEZfE95/LooyUKc1mZQQSEHTDY5VHkImJ1n
gTw2CyqAipO3R9xouLhtwU+Uwcb7Au/lpz0YTk8S2O80+7zsW1Kc+YNBZsm6RhWQBPZ9xvAObccv
9QR35pqpxLbg8ELgUfqKI53nR5RqO+tzcf1Pty5POizfmJq46cAdbwq3iNPfeD6M8Ck44A2LFdiV
SIpMkhQI53Qs0ItcdrhgsSzeOak9UYXx4YPEtdMdAgs0PS5i1pv8b/5yGCtuzRxxfCThFA5lmZnS
ZgvyOENnPu0PTK4Q6GYeg9IAmvrh4zxNfJ3SJWtNsjjYkRVr32Ci5BBTKjyyUBsq/Lj5x4OVv1rL
dw7Do206b/ZVkrulf93jz1g+ebG+JbgQ4akbsK9SdWsfaJZ5YiEU03rBPsSo/CIGPLV8tOIX9OWD
Nw/72IMAEQHqSB5LkJ5FxkHkfjpT3c+PZMAg+FfzqM7fWy+G3Eox8GIinqE0ZBl0VQzwg2j4Ge2v
QfEScUj301IW4uS6p5KSPXbHv0yM6SSzoqmtEk0V4q3Z1jxLYfiDf7S0+EFV7bcJfmosa+bR8Dqf
diF9XBC6EXcwNXVcaRqKbwwUv773z32xSC9i3TkVvMUCZrr/umMiFNyiBCuiVHkJL7qQEtx0T8zc
khV1jWcecMrj5F6gNSuxPo3OLEg4qeUsazDmhD2D/Cfbj4Ubd7JaMJT2oG3/XMpnbnPskX63MJg1
CBMfm58FjZsnJjVji/jYKfcId0/hzN444l6+/O1mu5a7oJJfx5PhDLKOg3IwIihkSKy19UIReiEz
igZYLpGh/koAtkjn5oaUaPYEx1dFwoOY7eYbUJ9o6jF5DRWMUTMdA+gVBCG13UCR2bZha+3S9VSJ
NWQdFxcxFt9kuHEjF0KJpMaTykCJ5exDy8o8Zkyuxwic1NK8I4gPRQ9FnoEvOjFRPgzX4v5bnEtB
uFDK/+WHkz9BpoZtWbd+s1HD8WAtdZ5lGyOOeNX19UmxI3Jvz+0KMj0LGy6nyXv4oUmFGv6QLhrt
FpSUveRzy9wejmtNzTYs4Xjx9VtLZsAQLIVvxXb31K37NiaDICdRlCXPf9YQMvK1I1XG37RlJ5fe
rAlPCiZBXycpL+VhguXGWlJ79jo0uZWJkha6y0Rzy2B35Fzuh3ibi/DFgCqD42EOUvaLZ4f7Q4xN
lvVxcgSsHyAtWwkg8kAj1ONFPaZWRIfeIaKnnFfwBVORmqwX4TLNOxb6QIAW2DNCdbo5NKSCO0w9
HkoxY7CAodPq5pUwhQUHrsIcos8TSQK3KpocS9bguCB4hWsc8/S8SlFFatIOZN9yNLZN15/qA2k+
obM927LsNaSi8tfEK6N/qPOLoFu9nrNXMmbtNFIYC4j7liAHouOpOkEwZmgWJpLdTz3c/tEN7ce8
U8M5tK+mLLytObzpsrOUdhklBDqo9p19j4q3NiKDtEqUTITdyBRtc8qQss83GWr29Qex9wsvH7V2
bw0tPO80Jp+fRVttLxVjl4gBF1I6mitPOnA5nGb6bSIg5tJ9DHMAYYHG7zY01naC76uA5IThSIuF
Dn0bBQWIf/OixbbiyKUirqGMtmUGBiF3QS9PNWeUA4yBpmbdPArkjY9gWcdLqbbJvTu+10jnGHHY
w8xwDj6hMjxhnhKXy87BdtwQ51GXLfLji3RUd/4cPB4XUsYITNoxinbCeXX03jI4zqqFNbY+5ry/
pxK7YDlg5GQEGwu2YnbSjUAuNqfGqXh5Pf4Gl5k5/IqoHt8e0FdNALmwaKwuMvs/lLLFmLMXcH7f
JN4sSq9y/t+Kh/r7gCGfMSKNDxuKfpAL1bpzeFCyuyoX7exoRCbEcaiBbGt/5vzpFyMBtvR++6j/
9lpME54f0TuBqVSfKLisYis3MoHgRcypgtBCDs9wlVpbfV6ieIytroOVyNm1vorGGeEziJCZ3S3/
htQa63Pn/zv6kXDQRYDPqj73mKEyIY+A128vbV7yzV1XHtNZrVksa7Y7XupWgmNFzgSQwHpOi6Xp
HQIvPIdR2+XXYVS6Wqoof7kviLHTdHj7Kp1pma3p3GfWxMedmCkghyuecR3+IzbImKZs/XLTybqo
0bRa1Z/CRzShh9Jn7QpWZkwKHo7XMCVPcp3IloTFgZbbz/obq0kmU7y03FUORvcGXDQ8f1qE/NUc
/DZ9um3LtvCaqB4qUtJ+WmTYjU0QzkzHf3veyfyFf2781a/7NqfPtMkjG1V/2cGTCzTkNKmfnw0r
o2Kc2FIUPaTtbIyO9xXOJrMw1XooSIRnqxcxf/LWcngZsP3WWEAEXU79Zf9o5JKGv0AeVO6wetl3
sMmoRY/uDJDHRMORLcfh8+yjRvHEXFO0/1ez/iv6hyeNw3lf5CjzlPChlDY8qzz6+A52KDqu3CxP
XgBhIDhUxavR+k+P/4aF3O/uIZGIU3UvCbG0t4w2R62gawu1PTH0tWAz6fISMGD4I/h+pcxc+jZM
z8XsLPID24aq3YbK1LbGaUq9R1n3ePGvKgIPh7/KApsb3Zpnw3cZ96S2YoMercYMlH9blx8DHHHW
53V2VVZyB5jSuWUcfeKsh+U2gxswP6MRg/dUjqKITSj8cZzhW+ARqv0ddHJcU+4k6LGOTZkvkhWH
JMo8Jc5BlcRekPovRkvEX4x0BMKXkf1wDnqb6pO4chpn/A3uP+kdJ75q1A38HTgyeAwop9T/TiR/
KHayEYPF73r2tKcdLvK0Sg6EUHUeV4mQF7yicjLIprrOPnqU/1rt5PggKcCpwIlFuk4ifA3m3vFI
jWBT9krfGH6T+iszle81CHklPvLEOLI26jbekryO5GSXW2iGLlyiGW4xrjpLLBpQtWtoqXOOiEyq
90+NwA0JvOUnKhcfBklc2lTwWRuF+kWtQ6eRrmGheQ8nRR3F545IZvGpM7Ljn/k93jjYGOdqEHbF
XM7horS1l7dhc5aknGL+zFQ89QkskxKTPmSKI8uRu8Y2rW/4OkU2Yq83tVTkGk1V3mmrLHz8JO7P
GnOTILSvrQoDgwPme+0RZNXdTpMp7y/k2ER6Mkug1k103ZeBX9Gm9BjP+nbyUk50T6sd6N/O1oJN
JElYSjnzbcpGp2RC2x62yLY10OkMYbTK8+OMCM2e3mRd5sxHwyPys1DVwbeudJCAgAw1xd1WLPSl
W3HsnFtlCgnOmfl8NlpUMfpWWwpAg2EVTBUxPvbv5KbQ5hEm5rxVqsVKgqj5c55udwbvO+GKaxMf
JEYnIlqtlpASlDwFyoGSutIXwwv8px2CshRImlK5ha+aFcDN8FRkwiM4gtsLdOH6g4p7JU+xXMj2
GYZQpwhCnCxjz7Dk1hIIxu3xVFQ32vjFZ0r6kBx8hNerh/u93P9cTnHQYbqOKhXSaxO+ovZcfjbH
BSNsM3A2KpwfiHWE0TyN/AdsgUSL/gXV/nWEbH2C4hri75KOx8whYnVCyq9XVUd1bIElVXlO0IrV
5p/cxoPT8RA6yuOvXe+nfY40GfaL+IFWwDln6qLGVIPulWb6iFPrrcZPkknAzmFyBBlscPk/hVd4
G2lyLfj1ZuxUnuLpHvogoR53379BrAI9z7rLxErp0A1Y7SfM2dUhEfRrAVhfw0SMh4Snw4mf+h/6
SbWSQCKQZBnbuSn8TbASR48WStbXZRQUfY9ZHAyBXLOt3Yap4DmUMtoQYvYCxRg3CNoREcUAvmuH
/Q64xnaEOlmOgrAAfNH4t1SJweKAN/2eiTznG6Qj98ab6VXBfcjSNcxSDc9yrvMeP+iRvnqqg2h3
1vwJzp3XQguAjJOaKTXazIGhAFBc8HMDjYu2lqBWUywOPcTUFMmAd63W01qJzOWFvQzsHkSFj/Xh
Hl1DqiwWkQax/lx5vhHybNKSljLVXeTlqjalmUwXOOYNhgtZNl8MJ7u0Y2jrfmTc4fIWbvTUdTxQ
CuLCUMXihuYOQLt6+I/aQVCHeTHOKKDjdpkjMU8Arwg2bO7FhIomKK7hvs5TiaaHfuF7jTBQAfKL
HFoZwTuF2kf9GOPoiVLLjKhxU/Wen1CrpwQWTfbOBfpV8lT3FxJLsokY36ESwv1aVrJG/Xh7gxUw
8La5fdTkXVVsAgyMMhMaJx71pCWjpzZ/qy/CnwBpdKbaNsUs/GWyo5njFFpvrQLcpaGqGfvGWOFv
HnLdKYDJAu33t+9xmgITMf9d8bY1FY/8SQ0ctzzn/LTjY52l0wxEyMRGfJAWa06Sruyrd5ira9Ew
n08HMEWsCDndYDISOQFZIrYAMjHakMzvLHYerDrHrHolL60OPkoZsCecaqf9gbodtrxiuDpHwITz
j5cDybtXU74NlsJTMcYYcyqyxoLst7LOmJYiDnZRJ+U5FYFuZeOY8gFJNcC7PpEw1YaU7xllnqpO
rc0RhfV0sNOk/une1fDCPDcQUUilJY1ugyOp+Akb1DL89xBYyuasvp+ccBvK5v40bopPxunMpiNN
QgyvqdDZtnPGTTvFxXmoXpLUbPRcLyPxcvAds7Dld9vxH+bglVeH55MYVRVy3YlybacQue/edaNv
RuiM5U3tIJBo6SecNpu1/BxE7dr/PyPihqwzIUdH7HzEbdjYc6Mil+OlqwP8yCD3vesvVw3rTXF2
EFw/8vA/ibxij4z6ctGFOqIdxISW2SVct041suj3rHqj4pbIepk7rnTIHAwDPuQsgkhKrnf5oQ8D
icUYiu3e68bNjPPWK2Pd9w/jJNpx4ZZ/xV0o297aAhkEr29G18ekxURG5Zc0LzelTMXEGBayNnKe
EfXWScS5m5UU5QSWoZGoxIe4diVmhOZMZ9xozFZClBIXGuAAVnOMiIpLFXtLpPY9PSCWvaUpalFu
qXMueSWKJRHvAZLpQ6e3OikhPF62kueVXSMC83aIGH/2emK3EFUNzEnoppsnI2r5GO6S68LjFcj3
Q0eb7JBx6py3x34LOKp2xMnC4pGkzqsLfqSZBLHjEt1OHb/eVIkLbVhqUzx/hhIBf7W7XbPvl988
2E0lcoNkjUYJ4WDRo5g0doKaM/D6gvaULpSgRDMsIRJQb0IvEXhUOszR3LETriFi7p7HaG20aoiw
PNy1NAqnOA6CqpdLOOgi8qU9PLJP8mvczXMtd4EPWDzcZz/n4JiifpuCmq4Bs7a8qOdTGHozeaq0
/4OoVavWZJGWBwwsXnIFwW58ZrQ9cg5Zvwtskm9cUtwgl88EnzCpcsUaSX1sMNp6M2HXLipd8IFX
KqgAW20frZBpeEqPx0WVEZPwTOZ6ba/K99wsoRYhBmsslbl5M0UiywWnpHrUf6HuF6thXb9eWPCj
PHPfLJ0Pmi3JA28kbLhT3RziPzVZ1M3HVHJ5cuI+REwfVqvJaEyLOWcT+9JbjL7xIQ7s5dNLK049
Iv0r4ZtTMkracB6+GWxIDintXr6FafKvvSlV9eesO7kX77fLIfvuGuNxoufKpzBSuA9SW8R2gOL+
449//PGojxJRSCYiysi82Fm+rZYehyV8YsQrvEzRcCfAMBX2/uph9CyTwx+gT+PZAe2Sx5KQQ/tY
vi+yz3WtqUSjPLM8PqRoE31TYDRnHg5U4Qe7cWhB+woyxdV7SRk1vByNezA3xjnVJBwvT5s2ODsg
IxgmrHont/D0QROHZsUyaPx3B3ccWAkrVh+NMt7rHgw74j6hTF8RgLsYYRP5pqdgtQuN02BtkagH
z8dfY9aOq12ZIqH4KftAHgLFas4mZlgvvh98Hnkh4O7OEogfMTC16X+vZm5tp2tAQrbewzccOBZC
nigwLnkJ92jGvE+3gTy1ALlRusck21spIOqbFmwot5anSJ44gyIQhqDqYPMVIl8Pg6V2er0GFcck
gESkKDpBskWazi6Rhys1gYHri+PdApPJynzxhahcTQRqXm96OrLH9c/8teyNNTVZoY5Fh3YeiQYm
PCylVqSATVExifHyhk04bb0V6Ska2se/XJJs4kqMbzdSVIUDrU0JQZAap6ZKyGDf4BE2THqBEXPv
YMsUxx3KoEJhQek1aykZqPZk+kl2O/SixzgVvT3hzX05Og2XQC+ev1yB8Pmwn3txg/YzkqYWDKjD
yO+v6g3wyAxnbBaIjBGZz4JGl9jnO6/2WnEvcTEong2z1N3D5MhRH+rWHdJeO1qOVSHvOL+5qQJf
MmNsYDrm1lzuig6h6ynKqzfAMSIg1o39ToXfxYukwnaxEvDxnzBg/QS23t6GLtLa6VhplU1xnzlx
N1VV3aWdCbHO7EdDvua0ClKNpE5SD8CRiXeVzUHa5Cu7yl3VDMnUs9XVtl+p3S0+6bj4jdZypx9I
4hsEGARguMs/mcWwa9WLl6c19H86j1pONiMK7YNjEjguGxGgdslxIIbCFcUKZvr2GP4SscgHryqj
0mGL89S5mzurxklW3q4YCSremNdeNVoziJG6VxAUIO4nW8+XVLEYkj2l9Auosmd6in1zZctXJ9bV
lXJuH1tw27Cp3dvbQyltgBBrHn9WCwBNMkWm4lGfyVb7eZfYzxOWYk92gIfWrHf11qVbAOFQcZwM
xnhOmhKtl97K922LHzOt+X2AKYdEBcMJ0+1Hd5XjDzaxj1iVYYsvMfjbpcRQQiQcScp8VvA/eW0U
zljN2zN6KUi/FD2GYoN0YLMcD+xe22D23vdfOdNnZMPdn1sYGfwY9VuFG51WrHhqeSObk2x0H27C
prvnVoA5Za0wSpmAPVzC3gs1TZflYRUjtdgaHRnc/daMfrDanO41GPDbXxXPohTd/0ZLu6vwUdic
ul6+prMjAjOvOg5okmWbBxU67chVhHVUZInVakAAMiW3d4yRMtzS0FRoeyiw1HJ9wWX3qMvfQ30U
otePiAkc8/5LoWAqW/PGsFmCNkyhAkgeFYNe27fFN+HP9rajgfmqMS7rM7yYmhEXr6qgLYLfLGSq
2yR7rUkUGakAid8eoWzDlbkIo46cK/RTTQoILBtRx95wIhfXUnugbEgHJSbG2+7mAGIy0UZqc5Dp
19J6fVU/g4KoARGyUoDUbfuFePxd9GxKlBRbdzg1uNDTDC/4Fcr792mTjNmcaIyuvdRokCCu9Xqo
BT9jFpoukjLgn2KeFd5TBqMJlp3ob2wR3LkbGPuxcRQ9v0wdGC6bGKbBFpBFxdeG6rn2tX+Qx+qt
sq5A7sHSmSLtZk2U7icYQ3PXJkkFORMq137Zfwx3UP1USJGNVSa9XA1IoscYdpJTIXPiC9+lNCdA
JOUbIoCs9zUMWpz1ZNwxhnbqQQ7AjpLL/X3XD3hySrJj1gJs73zoD8pxNxte/FxmxbNstejhPC4O
qWoWhg3x+Ce5QQOcFFPrl6XfVPpcy8HBu4rF4Z6a1eDfrXj4dZycVEfsbuKkip/YNgZ8E67+2zT3
PePPjDbxe6QGE9RCu0hF/UfkCHj1yPv2RPVgeHUvij+m3go/A+JU6jVY+eeu6Fi3m6zDTyo9v1ju
SGcoMNBMDv/gYQHXhpB1/DQyBUFmYSt3Wi1u8rKkmBJH6pNut65y47xpyc+1N7/x3JwyjVMfVH5u
3/YxYUKZoYqftuy378XanmxThf7S+eAZCyX/fU2ta6Os6Evd4AOFQQXc2Vn260o4ldcFLfLRax6V
vt/NL2bxUrhyBa/zYJWjmgiaH9nzKGl1ip+Y/XHpQIhqB2R81F1uRCUUr37KcPTTgBpD6pedFc5O
lVcB4HBvYAHqslYL5pXP3Rslaq8cX0M3jNqU8Z6B8MAW4SHPT060QFGrtDCfNG1iYfGcPC2RPATI
fbaCt/GbIGZVI33lhawNcDfTdnVcS1kvszZW8N2Zxb/08PiydzX+4hvn7PI6LMRnFR9aIBpWOBrM
vkgUf2cxGj+92FXdxCOwENlOHLjid+LOdGXei1NFy7Ussoe60GRsZsXWwr8pMoysQN/GsifraEGz
vts9WOKKf1qeKosgRX2i2tRgQ9GXmilXwdirl43EPzeZK+s2IhXs2vtSGpGKkNN6K+WjI2qQagP7
4hmdOXHMiz5yT7WWKBdf6DMnQC4klLoW/TBUJBU8JCFLUK4RF8hJgGG4/ViObj2aZxVBjjZUrnaF
ltfI/ihOP1cjWiSapL92+AT1+IazdlOiD/DrbRCej6o2oC1vfSXlPebjwhl04lHERfGKzYZtvvla
r09Y42JCYWLOTUQ47EdhG61+jVEnlwwVYLvYGmW15lfnXWmRyizJRozmN8E3YnRXze064yw8z653
4ZYd1ZLOYkUou+wdOMA+TeqsDN6OXYLpCQlQv213TcACtiY2ZwsSSFDTs21IvF6XBvyux+ynu+Tf
JqMygOTgcLSNoaDwNoMm4A8vp5fuOLD/JiabZ5DHgRyl+hVg/ZqhuuoOXGgOFWG09mQSeXxjOO3y
xjW7yz+PWxad4OAF8JkUU6U5J1Lf+SJVmf41PaYH/lBbDlzIu5tY6bihjqoCG2nSH95kfKaXe970
QLFDZsdmja6+igU49pkEzrExi5qzJrE3rr3q8C5OVzryl2DxCwC8dPHq9C+kWEpgQtDC+6GqJz1Y
BbOxi0iUoH4VR/ZdtgTYINsBUi8eMbCWczcFFi4jRZNAhf7P6bCakJK8pAu8BOSUAoaekTWyo5jb
yu+FEewvwpVCAxh5QllroZR05yYr0BBq7P3xTA7vvPT1puxkJckZQgr783XgcFewmV1aO2pWhshY
ZbNBav6nIrAyt+XmKmXK+3ptRCa+0xzEXEh2bzMJfjaMjkkMCNvSlFTn6tWHlfBA6gqa1tbr9BmB
wU/yGaYD94cCrU9VuTD5BD6qsZ5zJggGmRq0Bb0WmGCPnsIck/8jPSsvNURIJzllcOTQylJT43Wy
rACnnXOfRkRPAHUxDJSAspRUaBNL2H6fAhqlQxEd+6RZXnhNGIVHFZwyI4oY5TcIElz13mt1mjp2
IYhwEKYmWbrc9PRok2aRi5mYmFSHuf48+NPIAMnBI9ntREeQKTtTfKAfKH7JeHzOEiAL7b6B7drY
aqLRLCPnmXaTxN3xrj79U+jzEB8OPJjGKzpPeFMyw47+sMd7jclo2IVy3duL0hm8EMUmyST4nklR
MDw6N0yUC9xol3qIzIYISGhRKHofMtB7VQ2AmVIws9KXAd/aLp0cXNuiCSmuBJ0Tc3IOUDwNNv62
MtnC79XEpSqvF+EWZ8j9uL/geAdZHV6910kpL89H3Y4MpCfhdIoFFqLTlkoui3EkY2AfCxf+7izv
RJMf2NCS+bNY+tQpryLBr4tI7HnY32wtXlMdjmOJHbioSzUCVG14Cdsj+BkrTXuR+9pkeHkXn/J6
lTTAVFjZAy3FqfmSB10AyaZ45BHOulkmOa4Jb7RWOTqlmbYl5JnJy/4sGYUrzqS+Lepv8noXS2Wz
hRcd548Q3Xz4gDjd1k6OLYyTTkRuao/fIpX+D1s4jNm9BA1ZJEecD48rmAAyDiZ5jupX4NJ3Is3V
xzzEiCq5geUVaNM/WPyrfMm2br9RTtLs58iOSaXtWt4yr4U90Y393YRHQNS2WD1pjC9qViFJoBRZ
IP+diPI5pR9M3RXcLAfhypXwByPjAksrJ3bPcZ8Cb41xQBW4MK2JtgPN/seTI9frebcICmMQC3rN
F5y1PNWn9ggCijAHsRB1Z6XWsYlAh4vIrHQJEVTuSUdb5NsibUDANtaU9DZS8i8IR71vlEjm1yRm
i0vFsm7iZDcWdI/SbAK0tUILAbK2hL3IoM62esz0/6SwVsFpNgA8p4u1aO/2MSavDUlUNGxEpf6d
ECBY3pFpfE6q9xsHkANYoZ9Xq+61KTm1XGNspI5+Er0o0Vm6OY8YW99xHkZI/Tay9xWXz+X5PM0K
HzuMBGbDOUQ26f4gML7kXkydRtns1gKF5u0OeJdE6RHCobiyUn8MivNC694ZDlawVfqgfyeox8ot
OVOLerO+NrJV646EMdeCWd2G8LswD7K9Qt/DxN/rQOhViPsmvPvTkBlORh/8FzxZ3omGzPs1rsCp
34HYAHB6r06aizi/6HXoWp02MbPJjuBMWhx0O3nOAsAu7zr/OLnsCq5KZPSeu2U2MbS2o+1wpsqa
/G4gsm0CpdcSc360ba7qJHcE0oS1tdV2BNF1b8lcnfISB21ai7mcjt+qTLaVKycczQAPBxDLWcUY
rSRuZtqmXAMtZC67FSIOqcVR3udNtug/VRgrzFObUFD9MaNskcPbvfK5weKNlM7vZIriUfGEY/a5
WYnNFeTvKcTId1qNKv4TQs/DVztUobmtK3LAyLp/tSHx57mFY1WbuXyChRW8Oc37g1PXx2FkcmGA
Dc4sPutBDat7DvLVRBAWYhTRVYSRlTRqNsQXhLGMBoevYqA09K+REWvkyVr3kR3ACli8QnWEDJgo
y0aZvU6OzfGI45cnCj27O+ewJI5QGZ4Sq2QjIY2+CuehdrQ4hORYYZvSJRI2ZTQnxMWT2xZiZJXz
ygX7dWhgmny3M69yQVQQXkHOmp3gEc7wIL1U9Q9VzNcJPMg0KXrKToFtjbdX7xyVNBOntI5/NHqm
avGjqVWou2U8lYPfuJG7rQW8KYq5KQm4rRsQgeHhgdGsWPFLfLiHl5xAvHxkMMLNRdebR1dCTnLT
qno7AZLdRARfPKnrWE3uIfWqfmVWF9rBMSBVCydXjXz3B07yQ35FtnNfF62a4Y4RiAq3fna6z88N
MISFXeHWbEbhpre714g7jxVcpkSUf6YNQQUnWBu5k+yCm3OI8u5sEwob1shNpfTd2/fq5onaOa/O
MeCd8G1Pay+rQUN+tVbbqQZq+KzHC8l/CDAZHVUbBgRyEOkblwaZObgDWXGCI5sb0OFhttSxT2Nt
qpgrK5h6vOt2YGcjK62FoWDUJSFAKOk2Vu5JMxBdLYah7VlDg4bwKRNkdcuOWBwUh5AwCC3mWLiS
Be08UBotnn3kljwbTvQovbaOKLDmHJaYCxIZ7j9SjtUkX8nE7Y0VdVt0W3dePEEE+GqBunBgGdmK
IKrLt6h4UkpLyq2WvfSJB4JnWf9spPWL1Sf7YAEInOm/M/O7FHxoA62h4d0rH8nZHi9sqKI7PN2K
cKxHtVhvO4QEmkQ6y35SQWOnqgG3wlZlKef671PLUc0Z0tdOYFyvKuX9OW1pWu/aGvZRnQhN4+Gk
f59gwgqpsvtdlOGR1yxB2g9KiSSYS0/NGUJXAOwsUFYHBmakTijZ2eckoMDoJJaGTHOefX9Ym6LI
ZkK9rwxlEAYe5Dd76awsw7yC8KjPOwI1yQKnEvIO2Gp28Dwt2QKCk2lMN7PBIGXhb+nbWMCSz8+A
1mTaaKx80A4YYrK5uVr1DJWgaRZhuB8cSDCYKgMjXLZjWEnVa7QbuhLFBHKG0yMlCt11+tsssL8y
QKgS+JJR2o5b8vUSGK06y9IgqvGNHZ8l2xXRQI/rR4wfr+LqoJSd9U2QhwuO1WaG80X4GE6l3MMx
uE24zHjrEmz3PFJ13XnKqu5vknU3e7aQjJxsoGVqXpLLsc299Aotn5ay1hhFPigdCZwaZH2BucDN
fJNsKweIUF9IqNJ2ArvpqV+IhUoR9Wbk48lgg05GA/SrHfKRVF0T7wVThiOaRFeISeplub458D25
PW4Ee5sRCWbQOK66cIZRhj15IKhi/GDQTsDdc65kixs7akXGtNdiMSXm2tpG3V5yjv8BnPLogGvJ
UzGa3/pm7egTvypEI/FlcKJGLBXSInONqyrM0rt3vPO3dCWlCoLsb4I9JPJ4sMOfB3ZsyHPCvr9K
EWW628N0JZ6m5ZUdmAu06obkKnEx2b+BpXXjNPonBO9XW/QfGHoPvHkHDp2FvKxMVNOBQrWH+lfQ
8QMLCuF65B6JgPkD/YR9jqjCJnh72vxM3HmRg8oO7bXHx/K1mfYL/U0X96c5E4tEyfPqsLLb2+HP
9tBnMe56uDSYhy2HEq1g/f8ybRw8yRe/knG5pZ4msRq0c9kVIu5BV2TI1DojAp25WttAZvyIxMpT
Q5uluNb624oNAOH4QWjsq0zVNX5kWExZBqtqqZ1DNArnbntdeNv8oZGOvsiSfAnSt6LI84ZoGF6L
VublH6OJP89NjTFwgXk2pnTXj+qAjM98oDcFJCC2M+Y/0tK59STawfDlCn3aGDBurSa4ngCYF1Y/
GLx9EjjHz7KvqQ4ni64/IN7hJ6HUwQftG+HiFtobh1PrSnsb4ObwiddHcboRYA6dMUIk7/IQnWiY
anGnMug4R33ScnTRdVBkeCVKfTtqbsE8VDIk6zUliBRb/ryMRWYEveobOBJsSPQ/YQIv/I8jP7RC
zo601h6+xudlc8ojh+2WJFMp4zXSFIV1EwePMxseVIJDXg3eNx0+wCF2b7HBKBeB5TwNd+D95nyb
hXBRbh4Z10a95n4sd9iXc7uYlX7la1D/imHXD6fdyocByJ7PSotR1u0dS2OFiPCgA0C2rj8otBGI
ladOvKmlzBtNRPn9nCbWZ+qEifOcr5oxCvbathEYDL2bzFxCj11x9qxvleIyniGlpnLrbHfOZkPp
aosN2VwNrWsRcos1MDoHPpNBhbiLSKCzrgrOfiv7iX9BXRHXkAegrj1Dwj2MOBU1Tm3kFOb5q4xP
EMV3vWXpbn06HJKrL8Zr117djf0WYS8oNIVVwVGkeMN7Ia/2SWGVCfBr6oB+CAiaxLseORQst2oN
Zx1tYE919TRL1WvOg+QBqMewqxwwZvC3yfZT4U90jn5FcPSQ4GfOa+pqzNneKF/2LngIi610HH4H
8cCMofqsjyEwuIfW9CycazEJABexzbKUBFySoUHZXFxF4Z9djEQgS8AWx9YCdmL5TY7i6zJRxBd7
31FgkTVF9XwNULiMcQiMiS84Cpm6QXB2ZFFlnqqLf42IE8E4MoeGHJoLtQE7NiZBhlNDvqTDdRfm
JxWLS+yih0n+YNT3N7Oe88HItQH32uoMbll286PLrLZVquJeTRLccfBcRFylUjxK+/iGe5SbwddV
hUs7l2fJ6ZeMeaYanaLRDi2fWEhG7E6769QJYBEtHPPkMhoJwBFMRDDbNlvrq5qnx8pwfFoPhKJb
3PtV3yQkl07gDCMV9vc36VqxvzpcSQbXDz8zsuYLSJTPLR3zcO5VAB37wPiFYkMh5eGVvDDDL4KC
y16aKP7l5OC4XMQ8lXsknD8sEqjKegcgv/VywA2laa6YRVmjjwv2/gB+cuylYK33HEnTWDR8+wKW
rNZYt8wz6veIJ9l48DYTOzr5Ng4PsnvOwZ9BYHYlhkSBFNI0b7qW5XVtwfIxtS0kZCXXo/acACni
95uNHCe1K0Fu8ovq3zHCMe3Ebe84FxCmdvP9FGWBMN8Gb5XgjnzdPQG8+Tce9eiBsU4YK6yLOyEw
wjqZfw17fK6ZFkoJ0REnVFybKLFFojvrh0pvbrEPksbpNfHCxJmanFpj9NQDBJq3KpZyJxCyTq45
2nM+furXSps11ncOsdWDyGoIxjIftVoiDKI09E1kQDOYCBlRTzNR/zZ/3WEji0+ggyc56kB8v6e4
SvniJRIe04LlsQ74ECauLJaWbi2PMHo69DxDZUb8eM3lcEPToM1akcTnLWiy08MGlDoL/4e7zD5s
aO+GTSkR5EWkhONq1GGZMW+Crzt3XgFdMtnSzq3CrVsm2aNA+by3p1lenXA4d8dc4IxmZkabUivq
7gBUxnBfvBKXw4G9NanA5aetCXjKdS0GFr2qvScUkDffV8i/xKzKuBb+4NacDd3gqIhXvsHZsVGZ
3eo/xaCxBNHW+KxUWft9Jl5TyQeUo7SAmIQaimotCELVeVemeh+BWw0mB5Hu+AdjCmXkZPW/NV7y
IRj6ZXVohMtE7kjsEVPN7JXNG8ObC046gT8csLa0En2saGM0lp0KWfMSYnQDObMRO+q/MV97CdFY
HpOe1CbFiQGrkuev6cRb//tVu3dIBgOpknKdXA8h80TWr/Ax3y/8vk6djechJ9tbmtzExtNNTepG
Ui8hWdRUkpmuW47PC2FrFM8iCxlLLGsOBbfQZmNwMFDIOYNn+DgJdh0jqlJvuM41k1WJovKHT5Bv
zeYZD/E9wk6sYSEn3xQGeIXictBKH4cvz4QIPzGkBVVPqyuB2hFVpdkUqOdeoqEas6pFIp6khwxl
sWOmNpkI/hkvtZHexaU9ahacEuNhtWWC6Ym5LESQ/Sl9OCspUk4oX+PF86F7HQF/ZqFH2bgTzKSr
ReP+nex13UBBE+1z9RnU1M0JMOdqTymDSaEmGDJH7H2MpnarI3Xg5+YbSrB6jOnl5+TA2PprDUMo
CFDSUdwtnBIa63cwt+IAW6PGT4UtyV9sjLdO27FkRg/JbGyAXD5FNiIQw5VsrHjxdjRBHIjivgkb
PS+qTPTueF3SMoxoRO0oi4SroPxGvsA4QMpUPvpT4tJ8Sy6wkf4Lfoa3LxIgc2OlA5OMLZqi4QFP
sxvqyPxeQkQl3rhID+vrCZRvQ1exi12p+U5zx/9lNYL9L/C6ffrGhBlLQ7MJGI0NsASq9JoYt5lq
88zMzsW9RH2axkvJrxhqYCCN8HEd3eDNzLrh/LZJNvzXKmdxhoXz6CzSpVONbdze5wIVwMkEYlbw
0WFv+Z7T0CcyfwNPc0tpP+6quOaNSGBC10wJBsEvT/1FSXWikg3/PRbRAQctpegFNhj2rj9CqRYQ
DrCWyWhnGC41Q4hIN+kFSKNa9mP4zgQ29z0bBOwsj4trVNo4R76Ry96hJjGxuP99ee6KuM0sqrc/
NXjvdwkCzpNSR/gTfgCvC9svmcD/kt5qZh/ughITyRpTHo1lHFyIqcm6cvpOlgGhpJtL97KW+hPx
dUzw5yPGoLMNeZG/lOlNwM6ZEaqgYRly2TqOLgcFyigtr6ziNwR2GMP04lNRKZscAP2j8oEw5+4l
P+5hgoVmJLFFkZ5e47p6onxi0JZUa3XPaU0BeDGvntpnamc2qLHFWzXWlQoUAIDhKPgHj1xWeYKf
gZQ/reJv0hHGXvGPZD9ZoxsEwXRIEr+wxzf0d6Bo6D7IUiEntgSF/sdgjuEJI0EaOLYCu54SlvnT
YNV6mTHezLVLd6txiBu7UKTbUtzqLBzv9l+oR2K8di0j1oOfNIMFMLlB8rCqSZ51fOvA7jO6QxSM
F2kZVtnEo2HZW2fcvCyK+BJY1MEpgWjLcgHCDP734YZux+6xOOjAJE//dsvD+sbSf98cSNQXvKcA
sS2RrBkTlmTd3dBc1cS3zT3WpJbOCvi6DgjMb9HTcC0IGRc+yG0P49kVsFTEmr4jZVCDPLjzb09d
CHy1/ss/91BqsxeijtS5sDMRnvW/jbUCJ8nNFXS9Zj6hkZl7Yt5/Ohiv01GGz1Cw7cNjWBAObA47
8sTYnBHHD4oUJdb5DXwFU64P1YC3vjCJADXwnn5+MId1siTDMzVyD4Wbx6QGAlbO34eLAO9LQ91j
LWQpnXQnk/F5+XulDDW3c0QzqrqmSlOuzqzOQwcGzqDs+GHRBjUpx3mfjlTnYP6+fefO04B+F/xT
5cJVPBXjbhcX0viC0m43itjsMQ419BOwxbcP1D/mY7e+jCYOpZF2cJM+pH3w83mt7pwTtr46acLA
IzH7ln2i3KglCbxUG3+zqbJVCDrDxb2mGXDj3u0g5Q6aBX5Rl7kvEe9BmTEknIT9AsBfoQG6Kwsp
mNJn4sQJ7Gtx/CmchGsfywN+/Lkg0Q4f21jwLWSfrsL85cXhvv6g7UdeuIXPzdxNAn/NzbaXx3t3
Zk5Ipba2KEN4ZNrtbuiIGnVvdnYRS+QOTMqP5jctvp/SOQX143UBvHk/KpsSTuB38c+B9r2gI9ar
vra0MysBphnFjIjt0yMG8gZIevVXdS/QSUZOv4VJY1DjCt9VgPdM1fo32ZEQUpIG73usRd39khA6
XTEF7sbD8P2jXJqGsyTpK38FgEpRn1drRoaPwQC8ce4Ug1X9WXKHtcorLBZUtlIq42HTd2xVmFwD
W4Z7PKbqh4l3w8y1xdjbgOK2jH6EzSrn3GBpymVAj3Oq3y4g2bEYccY+y8CoSCm5WF8vQkA0z0pN
OV5G68urMeXbUfZ5p5EmrRtoGoRT1sZ1gKuA3hFyblb5Gi9un2owrbmdl44DtJYv8VnyTVG4Rh/C
PQhILLYBBVrW+oLBGiIxqqrHlW4o2X1RpEZs88065Wkxs68y6aq718XeWQFaSJEYOyfJ6LWclNRv
spGvJdAjJwkrFBh/yEmzShv7STv4iSeaP26jOKl5SQk68wsi6Rk4dW/uVl3+oIy6zC3CIPSv5iMX
CesgTosaGsNm3AK762XWP/6z16InhxLUZt7X2C0Erw/ZIRLMZYt1RE1/xpyl3P+TFlqgvc6V1X3g
4yI11SzZH7OlN80oSfu1YHkBD/HbSBCI+Q0cG8gvd/NPLUKfkJjn0YbUxXAFRwJQ4gkS/0sXaM65
G7PukJhuia/OD7uny91LbiGfpNgNKTjfQzgVstftB7xLsu1+LKHAc9LRtUJnRj7ad5MC7HcWOo/O
1tAS78n2g+xL2LbulRMMP/SYzNggtGf8oQdUCF5V2O2iANZMVg3ZqM3Jgeg9mOB8ArC80Jsb8zNp
hSEC5unDbJNcoqLy6tiaKpIgnRE2z8BOLMbAaMnho5HmC3Tsg1EeipayLjyp/eChTZwE4pY0ftA4
lYDc+lRJUWZRM4N20XWm1Pqhiu7hIlqm7twR7Qn1O83zTK3mXbnovL+B90WSOVdFr2E4VQPuXwcW
Ly1MXogXaJ7LIp3myePbXcAMO+Uv/yBux+9l05f5qQz/Ty6zJGNGgc0NX9lg91GThFBbCOhih6Xw
OLNJAOGmmbMhYyfSZR8zxyDKu3YFOTdYORjsEAyHl7FqYvBEptoAkS9SGdcrVdwXXmw6uLjSnez2
tk20MltzzxJX4Vyer8HGaWQDiNMz5hNYTy1xyrByGeLfCGAMGxTcRQudEIqOpJgqxhzyAFycoutX
eGtaFoZpf/y4VfDcGzP8TJLj3/TV5JxsZ72GQRKQWDYfbCHEdN/tlPwjK38Yjr0NPBfjqTAiX9GA
/P6g3g0gLBjiO+EUASMRiN+wYAZuE4gisJqlF2K77+IlgNn1L9qeWSiblRA0KNEXgK04qQt/NzEL
FuuUzo7x2x67txIl3j9xtXQy5iLBQEMEgbKSXXqzYC3hfQQ9gxkcKW8UGbRJiIXm0mno3EwZA15K
hQWG4vC1f1f/3SGOQI5+BcxnqgTfQcuzF+PPVWpkSTnShs5gzlAmKKTCrUx4jTlSWayEFnZKzmQR
m5GXkoRWRBC/TgQgBertsPTTKZwszfsDZ/e+92ux51mzsA4gQ1mAZh7wvhcL4Z186yFeeh6jvEEZ
WfVTa9ug2pqsJFrFrrLDi1FRKTB1koI+cZ6wDNNCaRg8bVwVEuTmu8S9sZ3SrJ3x8movEzqiyDru
AnVcJJfflaChPRkh7dyrxOTMS2PkEA8MDYm6Udt4VsbyMw0s3i8P69EJLtGkqfuMZk/V8FOM3w2H
qWhefPg/lh0RXnBVO1lE20+nCMUFSYjUU489thu9Z82j2845CBExX6h39OH9pPZFnB8YXjDPk1qt
ouzItHQhmB3s0HdyJTDDxbY7Y11bMMlA+xz1LGbe3NE5EvdGHU/Rdb+juxg4d7byuv5W1STKUefC
GU6Qh0CpK1fgGVgszNo6t9kkLNwsMHZ1dI8mu0s6NxT9Avg7jlg3B5Nx/S91XPl4V4LVHf1vDlqb
ydvUVbMGn9fnudWacoTgtjJwk1eXVhGRzVFeuERCijj4Mio6VxTX2K5FDqY6dolEekJxD3wXjpxd
gEJvRgxODp2TaUvRtqoDIAc1zNMB7lRcNmRS2iqsY4O0PxymM7hh8MiCcUNqYviFtzexK4/ulVlD
1N8Fv8LkVzaNqEBDWBpmSo0wI6bRj0RLZlIySphzAz5xbr858rN7jsTQ+jwNQXdW4QXqhToxzJeD
utepNUhYXRQ5Sq5rbm4oLoMpM4vchThv6cKKial7c8fKiDuUfm6xrf7XVXaT3Ga4VqyJybRdBJuq
QiL1iQCYqHRUjZxSNGQBoAqB32w1FiQ3gmJAow6XEsPpOOsHHHpxt6XcE2dAGhu9l6Sl5zGJhOf0
9pndcZLlmpfTrde/7m8ONQ5JyI2oE3yL9GUT6hfQqwJLHAPyq7BTNetRiFT8TMnveY0M24Ka03hg
h0EDRk2qjLfqDW99l1tJfuUSjXQWPt1ammqU1i6M118VtWDgGEQUkAWCLmLh2cAlP5XnzMWPJEXD
1cS/gYED0YduPRlW6ja1DIHkXPTwt6T7E/7v7Y3TxqIkmlUZ+6oBO/Nxg0Z1FZBD5c43gpKGdUeb
ruj9bYCFguyjCMnJtDp5u3Jrz3dkcAzVf7Q4BMbApXYXlZ29zeLoT3WcjgfmYa9gxUsoHB5K0O0T
ZEynGcjVBXw2Ja0HgJJb3V+aTIc+kPTd1/c7IANZC9ZJEj/+fxAy1Q0IXn47aaJl7OXy5oqey3SH
BoR3stfpJQgg+jLnLbZ5uatsQrx1XOJqdjzFjx1y1zdB6UkZc0mA8S/Myy0O3Ut0yqAwBMWx92yB
V3ug+8T8ZNDAN16yMxkjrq1nUEECCZqYAbEwajUOdYYH1zOWk29aXHCNaNZBEAuclhamGfgzCi7Q
x+U+GvzfcNVoqNyWTgnRB2xoHgYH5B+5l8OKZpKtjNarqatl7uDh1bN4jzyHV8ozXVK2e8dOSCv9
UqtmGKOu3vfeD0FoZAmJCt0eoZMbyMiBt9D7FjxJupBfzDRwaQl7xR/SIB9trvZ/2OVHiR8TJNsV
d3LM4D+LDVnVcgM1ZxQ/EjYu0ZunJqMCPNMf7E41mSp2PvKdMhayabh1JqkAIsHo1XJOJUigJwpb
6CSaSNEoFuqiR4w99NEW9hfpLWXoyRKliwW2lJVDBiXdJKD1NWGZZZ10bsnxHN+vKbuO5G1PHi5Z
kXjClsVdjeNjq/HUSrqf1mHEVGbcjmzdiT53hlo/j+N9fcSWMDKEwGaF2JOjeVW28VJh8sTm6s5+
MoBS4mbPqO+pXOEAX0OQEJ3AVHYe+0DIm2jews+CNVuaLWhNhkvnjNVpwyjz+QSc//6wyzu/rrhl
RcDxXxKlTe5VRuLaihp2P58KMERetxl4wOhhDHrQPImk4Cb301Hrv76uWnsOtxZ+9Bad7/R7jy3o
PZKHoGMmZrObbMKC5FMUG8Y+gzI7UhaypC7/XqxaoaSzXZ8Ub3V3Wr+CdrJFIg5phU9JDs0d9dHM
83yb8DYAizAYZPW3R+k2TNlK0tnRt1Pb/tlUbFOcp1xb9r2WMIaoa+S7wNgZHdt3s6SR7arsK/au
flT3WGpjZfVTfdml/F5sujv21h6CeZRVMtd3yrauTSeKs9mKhw18BweM0D7VUobadfxt3owZccbK
tLwrxkNtdn4TmLTDanRXuhp+uc/ZRpTFPJsgATqwTaeJvVslHDlE5q7KVB1TSJ++8zcAG/VXL7bt
0ykNIlRquea2QhURY3+g2iLCGEC4KYiRJMB02yC03qlW9nzIM17jwYexn9V5ZrttGgcSGO1NB39g
PaYbbuiz/A3a5tWEf15pfwFomQuqCWwjkK3IrszxaQLzL30PEN+CeT+i3aBW6Xj9P6yKtqLXCL12
BhsLYoKDumdillctwWrr96j/gmVN0SRQmZjoxqHyU2wdqDydJTLwL/uNX1/WULNUfuQZVScQN++A
srFWjwjzYmat1hF3Yqdis7L4MkKEZbP3CTU3jyiM+rgFZNE1YjCRWfUcYBl4E2L9T57VJo0mteFN
kVnfoHgsBj1WZ4D3YrkV1xJPDHCX9BrEnwEIERwPcn4kEGUuK5HYHWMBz0RYdvRpxqmx+g/Jmw1A
Ac9l9tJ8CLa4bRJ23L+sO+RAImRXmeLQc/+4uuazeNadlFfM3LEJfFqyjxLkiVbjen0wndRo8i6e
4vU1xn2aGH333F9bnnAmVr5hjPc2EJtlQvRiQolt8SENqWUkOVBNQmU+lZFM3XxKtbiTSENJHDoD
sUBjnXDo63n7/skXK350jhIHgHr/B2vR8mdFpot6fLnU93bM7HSPJijxrWY04+rfUeJ7GDnLYiuc
oZDfuJHrCchgQLzXHiEptRR0PAobLNdW48n4sWssYMnh3T63CgqDzlpsPr8ceQy9YMqM68ijII3i
rbm7EeTCaevV/08QiR863qTqk9HfR78ylHu1jmB5NvszbjJ1kvHZAHPZtYn7Nyuf/4PtcLGXBsIA
PgXuazjUO574+BUd1FYxIFd4Gf7RaX5ItPvbbUsSrOMHyu4BYH+xZxZccB8sLdt+21QX0MOE2hOR
C5yd+YQdm1Ye5rdrNWdkaewhRHgGt7tOzNiyU+seccGKfyL0CQWSG9WriOiIdI3rthZdtCXl07n1
Ekch2KpXoR9CLQIAKv01D5HwsRJI7hFkTA8aGl5DfIIHVOmw85B1FLBJ4vQV1AkGt4NI70t6U+/k
Pu8bKwrF/55CCaBk/Ty2B+M7uweMRfQpBhJkB22+f0bHlt8hnjO42UC64064jS6bh94DSvVW4FkQ
Yv1e/tsntI02GOvvsegmyosB9pb6BuFBrEZeJ6pWPM+9MqJUIJU0hdyH3I9Ig6vQqUYGU018kycD
zfSzZMGJcwofzV8lHAW8KOBJur0L004QTN6dROTCoMrL282h35l+q7sB02377Gb8yM+BuXZ8MSVd
NMFMYr3N2Mxwk7MdsiPsaof9echqk9L9zLd8wZwp/18AuPFIcjN+hJ/tX2QKv/wjmZWOpfKYnUsD
H4VYq2jFBeOXhI0gxFUKo61VLOEixYVTXvGkzgBE4GjICPJ1AvstkzAnQJoJeqyE7aRBCiacJBjX
PokcuUurVEdk8wrP611fp8hGHrQo8vq9mTA/tBJcP7PZ9BMwgQv8CXVtRkc0oVSGw+8pyy5b75RZ
T5lAtFmg9HvJ4J1NRpG9iao+9gv/RDKDfjo2OvXcn8EZI+HCwLfrI9RywzloZuvEWw+0QTCJJxVi
Z/+9845OcZdpf+PzS9RrcesGPeFyWiw5aZIeYWzKC8RzLbTGAFMlvh3ZayJVR99khSK5BuudOkaC
lMZtqqM5a/LEfE67kOsUPtvMcI2seOk4de8QYHD0u/ychFsljNJ0bvcZelvXC2cgdbu9JZDtiDaw
g+YXlHaqBOEO1QnXH951wh6A7kENuo0w6bTjelWNUGlJ9C11y9eUbic6yjD2boFinH8cKnl6LDDa
H8JgZISfBVDPRj/0gSxZUytSNxInnqlhQ3OBUF9/QLBnAutLjl4VyHrjEGZSZCw/vUefU9HPeq03
jGhj3k1TsVcdQB1twh2UVI89WLG3YdhU57MYE7yU/gXmFWRAoRk0t6oyDt7SG8ca1WmIzov8a/21
cjGXMjK53fbQGkg25LAxpIZtO7Wy3mnxhoCZoO9aBGaP1d14Hu6y8qgTd3CSP139TJghDBBoNUxZ
RVAE20b10s0oas36T1LnnBU2356JogZ49e4EDwTvH8YOfafaWGJ7RY+l3veiZvEqydyiyqswrTR8
fbDX05aIPV9zFx7sSPefp3fmDdt4pUSO2m9pAtQDvD57KGKpgnp1t7gwuf+rinF1PgPtQh9/mDBm
Os2IBCnLYacGEk2X3WpT0mKG/WSdRvjbeiBYy2Y1Z03WtNzyMZeL7wx7MJxAeQUqVt+QoFlQBszX
BjuaUPdgV+tZHGwAHcrX8gzum4F/RM9sNNSo6F9mFTls/kBTK87KJwfpqtUc+3jFpCB4ggj8MQcR
mPy6gWsCo3Fnq6Y9GRjWe+DQyfNQKl07AWfQGRponlpuyJgkWOIw+BoHFNypgxdl4FfRBU5hPuwz
X0Y3Jswh25dAVZsff9nqJd6cA2BOZVPX+CWGBTMrLDXzT2XNHwneqU23y/yt/ySKnDq+735FoPuB
NvO2ncGGMwTp6sQCb3htqtFkn9tyAZaLhKi/iX2kOK6lYige6RdLGk1oriE2Msv3WtMDDRmEPS+J
Nyvx3hxiXRJrBBZr8veLszH35Y12mHb06i4F0YjyeXEY7jnDmgreYFnbWaEY7OO+af65KBq2kh5a
LX35+Ik9UvW8VE3lFdCmJ+U/kIF5YRS2Hd6JNVLdPoV2iEvCnCQnjy4N7rVlLrS9YK19yQ+0lBzZ
/l3KvMJJiFyBRyFO0S+SU3Qu67yx7ENb9bevDlU1N+rdsOYXsFDTFxqe5OYJBzkLC4NdkwzkuI/O
AxXgjMUzvsFZ543mYUZISDlNHApbg08e1l18IX3/CyLrERcHyUaNai9cJ+dAMfyR4Bg++ribLaHs
8JhacnJDm11U9/Ig9J6YTt419naiWaxG7BcTRZY0W1B3KZvTDWSljXBE/eGPytfYb9rDBG37Vz68
ohj/OuEHjZr8wX5STWG72MAHQsrBMKMM++D2LbBZH+JUlCqU/1+Bx2dVaONaiw8ZFOI6a9GStjeJ
UJgGd/pygLMCRVKlW8xmiHi/umir2BwdcZnniWCXgZLwwVrhg8WvaFV16PZMVynqm8hJ/VAsFTH6
tllzy/FXGKa4vntH7JjrWsGMw1Qi+e0rI3LVRKrQl9UsCFTfWD8CUhZ4uoK1iiBgPoM/y4aecDm2
6Oq7mItJuHBGhX8x50hEGlXLjFgBX0yUF2JCojGoXe+F9inB6TddDJmcxsgZChwt+PnbgXk3W24t
228m+iKfEjUNnuc1RrIWVdeWqUlkMtwbo/fRbP3ro9FWQE6DpLpfusZA+uoeH78eT66s0FKFoI3+
mclX561DUKkLq7Wt/gP+4TpH7VES49K5IFcX2TMCCMAmQZ2Yg5GKLp5HoR1IBwA+fDl19CrR4VSw
N/fEFnwGk0fhEXQX7R7yiCXiMTS1c34vF4w54XfgbUquj1d2NKIqA+2AW1IjVYuwqDJUFixAvvlD
xUhLRwCT/FNg4GynxRBx/mV7YRSptoBNBkCsx+S7guMusrDXt6/XjiKRd3gkktafJmuaMaOmEMPD
oqmnv4jMr2aSWrnBrgiKqAUaOS4wcpAVf/b5Yft6av3PxEQ0ZTROObuHI5q74vmy/6npUybpwmEK
6FbFFGDvkkEp2+OLfll6AUiHe2U6xOkTRopk479hszZ37SBc4wyMtYsdsJ2uXcjFZzjCEveEQVzN
tuZdF4T/gZkHbW6nkZUTLv9Fxorr2OpDMyavOBFIli9fPepu96uTI8Qj8t3yfnl1Il2pFNbixQK+
F4tWHPZDvhDhG5rEU08H989quXjUWUTtxUlw3V7hEK1D/FI+YRQ6YBPcDjDbxla+oQDZIiEiSYzF
+Ndg0F0GGT/7xJTm5UxVEEXTFxSnzpRPNAki0Dk10ZZYkRGKWC7eWACGL0cfTmFxOoloP8zgGG8z
+OvUWWAauDabdRvAa/900EnX8hQvwxAMeikhMOAKRZVikJooW0j8LwXqc2cmGGZXai8UYBRZWXgr
jhDGvuIXbAOj2EznyfaQmpGiFze78vFQn6agiCFP7It4kqG85xjjwAbYr34PIxBTp7Xdib0NzdRc
vGomDeDsc6aHeag3IWg3FSFXREg6HB3ZogSG+jYo35u9fbMEB2TMtYgNIxgyJ7vIINUe54ShHBtt
ezU725+9nSoGyBYvUMTKcvvUtfiq74WYW56H+IKIVylPXB4kKRZydAetMDSMtumB6EAEKAF5FBTI
wnxfron8/LeHUmM94pZj55XWC8ABYfasEndYUIPGhhYTtJOo9ySOSs70gStmN5WyD/jn8wqNChgR
rVQ23AgUCOdVPeb5BhV2PMRY8zPGD48XZ+/6q2oTGf4Xjch2o6MAreugWhdoHmoIQ3dd7dHaZpI9
2D3EZaPuztErVP+dUwFNsv9RYlV28/jC42BoaGQuLWSkaYl8Uh4jmDSnEh2uWMX/6Cw39AIT/e4H
FRlZ6XSEs9mFFt5c6Hy+6tbTJXN8X2gv0RbiY4V6uDNHRljRgw7vv0zE83fmFDkPtFBPdzex/sqB
n1ZwKMXxeMr3dsfYav9x01e/AonqR4TawLgCD5AJoN+8qFCaPdg6o0DmLjNzsE1jLbsA6j6cAzxR
e6kxOTb4U2R1iEhFRFUlJkkle6k4ZNHHC5WTckz3X/EP89cPia5O0WlRmA0TosWtCwOMtXy0USSc
l+LS0kO5D2qCM+QD8/pl5dDGkeqJVqXCFuHIkPlSpXecUDPxrPuiQcml9CWHRvx8dZ0SoUjcdJjy
Eq/FV7KGhNIKm3090dUFJB8XbZ7eyqEDd8DdpCF6WDpSYR2BpoFzsGxIvv0EQYvgkL0MLgSzrNg8
lh7OQEQtDp4iMSx3v3hz37sUJE4ZQYsag6rvST06oCUDRvi26MkHhJwVpSfxuYaHu6c3NrmNhyfG
KC5xnEs7PYHhPqpz8/YFvVuQA8PcFLDAkf1OLAPqB/bfBuX5dr53x1K7ny2FSKKIdxw59V+ZZio6
b3EvtTBAqW3d8eUyg5XT1wFY/K4NADQyMXvGnVJVlfFgFfdEn/w+QblQb3xUaTamin9j8S/88H4l
+0gaCHPyCisQSnA1lPIYeTdYWnhRSc/nVfHF7ODLBs8ReMqAgniS5a9BlMHGU1NLAcHku9l+km7E
BAvFt07HRAKmLxQQWAkDsxKHmRE1eXE8weeXmF9dNi6ktNiY/9bsziUAhHQaV415HJdF5M4s49G/
lCSD8W5ytevNDbPTHgjKhbxlYi8NsiPAAeM/VyG7TpE4A1QboMeZfuR0A9t4AyV4jMsaI8QqHuUV
XPnd6gbClmGUFeqL3ysQuV2AJGju2QvYozVSdhjTxaiWi0SokNOklG9ZnJKWr02btePodX8rg8oS
7pbxQ+KhpwsY8t71vd77AJWWctu5kw4ozXgitfyViYc4TivWiY6v2K1M2ZOP428xKKExkkBd49UA
+bj8uHxn6XWsYlMhWL+tmsidJTVsiJXVd9S1ec3bMseeZ9Bm+Dcn3pwnZ5L41ODqvLQssvM5Ia9/
zMu4e/nfhdVurojZvXSwpEfqA+aBkMsPpUf0r85fW50X7BNemHBAHtez2bG4wmJscPnp1nm15LAU
+Lw/pbkwZP29sJeIdsXuYDbkE8v5rK9DqxsJfifC0agcBL6xN/HJga2koI9xJQ/qT+qqytGp1M3R
MxtHRlypcvN1ghCHJqpEcyarF8kkZEcXZ3YORxgbQWTTvrW4K6IwdanE1T4WBgDemwrRQLnPtedw
9ysY6yO3grUqX52ndz/RflwTDJ+6Z+9DQppT1rUgKi8dzCQjKuV/DTCiNG5YiopI+30IJSTZhtva
a3RVLmP/ZltKHtx3aPLhRQKRhXWETw0ZxZ/837lDeMqXsd1Rf2SQkOPguhngryymBSKHjoNCpQF1
IIn6GIebXXxCYMvDYMtWOqqRoKDjPth5pZlLl0mCHr7jxbkA3fGn7SH1rOOJcYccKPq/rtxKAjP2
lPmVWPWJ5CkjWJEXyKjeii4Wlc1egb1GwVwR9vYFzyZPM1HyKhEvmzufE13UGz/CT5/s0FhWl2sw
gFUKPGHtkz3y7hpbzpQIfnbWPBd+N5KgrP2ELIx3uOdGMbLyGU5vUjAOtjztOeHUD9ZWZUCcOBt+
cwvDcwx33ex0RH4sWQA/405qsYyt+umWAKXtszkYkLUiyOBtpmj1fBHatiSvd9e9dmYvYO2KkGJk
1CZ142dnps9+doQbqlfsE7R/ip3JMVWdRUk9laFCyThf3t5R+U+6Kg/yt1qjUm2nubAkqtNOXA66
xGx0ryOWseAg692TJOg2szI9IWxH6LqNecftZaTO5pERlUVOVNL6FoPboOGOD9jVLXBxUWjDTg8f
Ixfx6NCe1KZ87vXus/rCKf+Hfi+/Px/rG7yPXZSNzJwTuKDvf5dqldz5+XUtmFkQq4JeQ61fh3hu
7ebqY7pm9i1+BJUMhUplGCY66pNNYAaGqWrNTpRZjMlETU2JayoYZdNZS5/nIffR4qTkEJY0zYqU
m58y7RXCiq7XbPXJDFRErx7I5CevAvo6wFP7X/bgiiBzCNxgwWIKdiPidVYciZdQBxdMyvHD2lBG
o1GeJsgaQqw3+vtlwbQzUsD7YOYCaCqoU/dvgSAlZU1P34S5MEIYOY25LD6rilzuJoE5vAC51gIE
6jqmNMfRhYPF8u9IeR7YjOElZziK3LegEjQ9kzMXefflK0lPRevAXaXCmrCkaHTJrSxwDR1/IaDM
ObR5qbHWF+3i/X5FNfGyQ/W/+lnqNyTmeudBFp5vgvMyq4HzpRizX8jgIsPUTQZhUxmea3MNijbT
jaaWVsfNwfwcX3lHES+TFqHt1q2tNoP7uNXQYH815I7O2VLNPL0+coQcs3toMvI4arR4bgnEEQKy
Bfb0b2TGWFIkpA+KptPvvuSvaycDLGQchkHI3DyOn5h5ZAla0JMa45uSZIetjgWfKtlmJD2PaNjk
LnSqewf+ArrLc2Dr4h8rJ/M9QVbr4CPKuBzvm3TtNUfbd9ilRCNHKp9KYQ6XLLZvjCKayfx1IPz4
Vh9ind9QLM7+w/iElGvRkHpOGQD/yhsaHOk0q+Cwl+tfKt+TLNopDe0/Kx3hw9bZbeBt/rDWLoyR
9yMa/0OZE1CV0Pk9Y/ES69MiCin+K3cL5AiAEU5Guq951jhKe7WhG5aEcEGmbMNz/zCp3rsf3ZH+
kT/nSuBnwxe3P2fK6Nx8F9/20YOupz4PVwUGtGrKIO36OAOi3ySxl7Ta3wmy0WTDprY41YBRDcJN
Gvj7dmKV8h3W6fztN3YFyQMc2mE/iY93D5vYKzlHdiI0dHR9Vbl3pzRMwv3Sl2hsf47j9ptg27H/
6r6cFG+P/oSNxQT4BciwVyjPG5V/SBW2Jym/TTfh0bb9Y5KM7dyWqffoYV9GybvyCPnciV8njUWq
mk/lIR/qKiEUuAQGvdaFYLKo3qBDhslKejEeoEJwU/413q5z7uHOhOFilvMddi8cAiU2l24rOEUP
LyYNU1r7cNBZei9mkl9N6eZxfmZNoa1p3Mg3XWOjTIALESEc6VY5VSjQLrJ9HAsSemvQkpGEImyv
xUmJfyYWX63dyXpUp1u55/rFUFCbPnuBK1l4WQv6e7U5xA2S1Lwi5+OUWFeZZs+wZPwfF0W0z0Gd
qaFHWHWgSb2ZBMEGhRmAdfNNjwlXRDGdTeHhY1Hy0bGX2ybH61CwIrTFWmXf7PgtVWVYVse+siw4
Vxa59PL9giBy2ctw+206M7seBLP6K+iavXvznX3PnttrBiOAI9Mqc2lp9pLkCWzeIB7DSja09ks5
rh6rW4BFJpRjNbJNmy/ho36p+M+hzxKS3QXFJz/T34yRgvk0BXsxn0CcXsq3iwoQTc5BatYS//Zr
SdnBtxu5MMmN6X252y/DQ5HfQLHQqwmvjaLA3tgYQ1FGtk33+mW2fIkyu1z7E7kzjaIhqinN25tJ
mCJyLzK12Qjc/UT7i5YosaDU/+W5teTMRMKchHQQsLvnu0Sou31KXHuSdsyMvMKHLznGtAjzixtt
CDG+7TK31ic/JWMXWgsxWuCXUdTOo54ghGsCcqK1QthpTesuf4Rqj2xwbWNCvBSSqHHnIAaPNbqr
8mXDJN9ekbbDfCt5x+vg0kND0+iBSQivcyC+3OirZlMfTcHnW6UvI6KRi/CdJuTjYkqqmXDHVYY+
0Zdz+b4gs1dwpF/PiH8A6FXGXOZUlEMOoeLjR1/TAmGK5zRAs9hyd3VbdDktfJwKrVZbXzU5Od+q
Un/77HThQSKtxm2xlYvW/HA6yg5a31BVFb1c0+N0JTa8C3rS5OWHm+D8yUmuLCnRU4mUCuKs9hGV
r0543IHioHxhuE7EUCQ5YmD2r6Jb6pw6jG9f5V1KhhW1pNodjOJzugh45/N5Ykbk58GGgLTdMUhU
yu5Dys4XmlLm6tNsWvf6OsKvxKpKsQuIRIE/uw/YnFwhbVg79Nr9RbJ9k8NoWL63ll8+Vgf9MQcQ
TLo4fIJoMuFdcVrMAvzjRUXWibrMZm5edvh3PRif8BDl8nKCXJT8SbtVEn30ws7uj4ZpHOfAdxHL
TzQDZrhDUf9ZB6WIqQIHCJ+z+Bxd+UUi/gOiLzuK+QZirrh9JOuNWCottEteeZe1AUE+rL9nbTva
Q67KOuLH0f6jy0uUgzpQgdc4z0NBHgv3mqszNB50W9TpBCYzydrA637IJPgol4hq2PMoYxF3RbQb
dcJ3ybuf0+WQ58OAYLYmjCPS9LJpi5Nf7c5Bp3Jq1PGpnzSF5rIYurl4Uep/1RsXj8gEtT9k/dhC
xJ6ko2kmDvgvZGqncN1LjdVH/HXmX5dSdvfrpF7g+h/BwuxSEapoUDDqrYHrXe/Taxy11UbxeEHC
2TrORvX4YOzYlUsMN5Zq/fV0svWGD/UXmGxTOld+ErJ5HC/M5jRyiqGsqZt/dNzffaHIbA0S9ba2
0yKXsklrc8LY8MGrLe19RKwodV8QQ72oOJJOtJujQh+Kpk9yq8knAh/2K89PMa0WrD7CmmWGJpWO
rDcSV2FrcjUTwWcP5dF1S07u1ThDX81DMEvbw860ikx+r3AoeDjh8yKtLWWs97PeG1CV6nVxN6Qp
sB837ZKw26hnIAdnDuFxJTMzCBmzn07LSh8VfWIvTsN7kDNp295cqBIMiiAnEYTMMmT656qW0WX4
QqUP3MO28aM+zSZ9wbD73B3ELsEXxgv0sowEQ8QubNbVyIHo5LcRn6m8QJt5h4N9ClB4s0DYG90x
oJQS7IOlTySH14t5SzyFfkn2KDLqCKkNndzU1woEQZW3QNdr9pVvGYQgBsnf+s/5KjdL3NBCyalE
4NaQVh/fgPjCbkON9NqOXYNYzHN7tka4tVWU8VlsBGCeM0qfb+lBaaHyaAMIHkLqpOhtuKW6y4l6
P+C9lyQ9JjEDqn5ra88Anay9eZappRp2EJi8tDNjhVFeO2w6BamoT5M2zy+liKjDS1JxeDSipAhM
Pzl2sq8Uv6LA3C8ogjadnrdKkMk0Y01UncMLFYZxQhavTxrIb99NIPn9yNNNAa8t+Zi1xLB1MZ2W
sOlaR04CbEXQDNqM4TZAyBvSbpR3J4rqFkUyugKc2AhX28RNMpiAMlgyN0PD+8Afor0iF4NWCUZh
WGauSwjcc8fMvv9+vVk9zV/acJ9zF2n+XimvfsQB2z0dKa7PMUwa663tefSTbQ3RvgXoXGxPUUeA
KunQ9sT9H5psWkRSQQuf4/8qj9d4YVTLgT9YTYOAl1Iu4ygCFOzw50NZPR8tzCTwLH999QCTfYyG
FDWkPJ6PJAAsogrcpKNCOXETsx17YL40VkU7FEtV6NoCWJ8H6ZYMPDTu81cxMCuqlPMI9M+afNHV
77s/u2UTK5//bAbc/fraSGDiAAA0xwHZ6J0AWl8L2L0RZHmuxHtiKu3LFt4M+F4fPvMzGnq0KU7s
M8VfxVUZ4WumkqgqtJnEeNDU7acHKQmMgWfMKI3sbAraYBZAciYCb9AeB4S5pWeL9UArA5Qf34rx
qW58pg3xWqLPJgAqA797ADJqwph5jN9hlGnqRskQPOhaxgIEmvkwLIAYBUh5YZH780kMtr9ou/LI
aunsot7JFD2wqBxYCi3IggcvvRyAvT1HP2eJb8WPleCRSA1tX9SfL7nHxa5aNBo6ezOWoC94IvrC
H01z2/lVJ32IARFkdybX7l0Jr7hjyHZtNkYGqgKRVCj8ph6SD+SQu26ZtCyAsgEr8F5eYL3NIy8B
K5SdunTMgFO9igr3NAyUKKQOJtl6cpmmjG96PH3Mg/KTv+yKsPpjtVfcx7JOPumpagT/qCEgt17K
4Db7v3it5kaRVO6wT/PSjAGGx3y+5ZlXWP+lwh0bHhaQLleQ3oeHKgJRQ1/UsOJ0NMHHNKtyoYVc
fPmheH1wo+GN824w/vqR3AxJSMPHbabHU7ajGbyjLpkVHDCRvtlaLqsSSu6j+ozKM78GgLe7muys
nlDbH67PIB1xkJQ4MiJsGFNZrT3pMCzf+BFjiTCnNxzcdu2fRAKIBM0Q0WEthoDXtttJc7pp0xY4
oAbDxeO847UERNagfXivFjPcvuftlc/35Zob5YuvXID+4Qx3UxuqwAV+Q9MaxYmHjKGoO0tay4lQ
e60FWCpehaqNo1VcxBl83FQb4XEDofQnz6k9ZglFBj2PJD0Txi9HeQSHH4tlbEXRofByYsleP84+
qh6aTZ+mmoBOQhsijrXADdLTqpMxsGLH/6t9qyip/tiexyuSOSmtXVGbl1pze0Jc4/axc2BkV40A
QC2uUUFIgpYbz8KFwp6k2IlCkGQA+KGs24AiuBU/7ZOFz8iK9UxlWDGH4Ur4GCSvYHjul/090x79
AuF872P7ClwA3kR0fpj8J0drN0P0JXqtHN9CO7bhHESMtg+k21giGcKTM9OLtHpxiSaDotkzhaFh
VKg+vIStmWOBJNEd1vNqy65Ty4mW0CR+SsgoZZoN0lgSJ3jhuLKkdX99Ga3ZokfWH+CVY4t+Dm4n
xabETRflU2NZVYVYJ0r+Y8nlEUEMiBJki7cIEe7K9S1tIRpxdhvwEGHBRZJyENk2X23QaG7aHzK4
kSiUZWlY4pAsp8h0qhqdcEyGi5p6WYynk1SBSGKlJosrJNdCwC/w6WvbTUUlp63+JdVtdAkvc/1n
bw8YsHLIlTuTNaSdp8uAY03kRTm/x71cZv3LJh4ZTZVi4rogOGnjWUlY4LIBPXJ/JPWAuNmQT7XE
tdZEbfjizRFNMoSt6UJ0JiQOajhnFT04nYkvN7jCwyJr4mw7y+mEvu0S2zVaJyyf1QDbE8GMPEuU
xSQJC0vE15TVG2VvjoC3jeyjzxhDZ2sdq5wSKHZTWcnAwU793hHdZSAcHinBdBJA0ZUB3XAAObAW
16HkFpJwmwOqdo47ZDqDd3xVitC7fojqsmoRQIYIuspiKSscK4VxnWkw4sKfF+6Ncd1rcTRB7fIK
prAzsOREArVfOUYTRR9cR+ZlV7aFOlQ+wmJ4+w1/izlzeIg4x4uBQ4KahHdXKQlaUYzq31+r4xy1
VOROZGdfpvfmaVPtm//1O4DQxq2QD+fbq/mB9IQYpTsifoCaB//1opBUcyjVnEnBUbddiq39gmmf
1pnK+SF5H8zNNKPzOrS9mZgCIF2M72fgvaawW134HdKc16BEAn2dnQHOyZHLOsKStpGSzWhOtxrp
doZirOZsEwOyskTv8J6nLpYlfqoA1Cge+mjaPM+iq4QrnmjgThnsLPO+GKVTSutDWtsy4S/jASWg
DCWVkFDKxm+VaQirwoJiu1aQJMpl9p2TRlzaRCg7sxdgX3cEakgDIZmn2ZheTmkfDKfL8TfCdGUF
jZzHdCHPxaKn9Gy2kLEp8r8P/AA/4mwlWDCeD8k6mQzw6KPqbA451FtnpB+BtDyJASX7WGyr8rzK
Xjz2zFGWpVLQevebmY8VsXbolAEYI0bxIwBkKt69dkQXY6IrPz6nuWrTVlRxU4Jm7gAgKnXlTc6W
sB7MpewP/h7LivjowSWBmcfhB/WMK0iEsIedQKo/O7+tY5y0NDzrjx2ZMtELP7JnbgnOnugq6voa
1QzKSd4KC2qqcUniAc7/FNcmnGaz5PecWArbSNMo86s5qBAO2G31vPkc6BQ4fUEybsRWdGdc66bd
jiGnxVnd5SAleIOU8UNzxaQ889e3n8mkoGcnbuS5f/MrRiZqz+IFx+3Tv/RrXkK8iiZQZ7DvbpHY
2Lr0648Sqee9SmBkTjF5mQ5vkubb9z9N+OQf93Sw5ck655aR1DZaMZFKdnuaPs6bhJ9El4botyQs
8cliVPLluR/PD68uNdR6tTKBXDGNvsAuaA4/Xd+0WI+lxhpnYaB/hZwsPW31YX+tWfOwNKHYXfE4
G2q6WBts3qY7ECc0ERofLwGtPj7In8uV+/ucDAIBwURUQ2n/D+plq8KI4x9d5o3QnuC6F4Xz16d4
6ztUkD2/RQLPCY9aoOlPi/qSmhtVimWjaE0XH3q9ODzi40yw+ntgfdT3TtKhcYF4/gdCMee1bJBV
XtmBAF6cR5ZVRq9PeKn25JK7oI2AWVKiZlhM4UC1A4dWJd3gQA2YjgAoRK2EExkIjWtfayKoAg+v
Ei8qtPfHcL9jxzzKXAA6qqRsP8L/pFdwaPe1DOFDo3Pwkmrd/zR8aSGysZqdgv3I6Or2Ca/DTZ9z
3dz9rQxXNm7LHnz6CXMzmPEflaH3it9Yk7IAXKGqkEy14g2oIf9yVRd5A87UdRCowfjqtGgJk0Um
oCDiwmSPq5uEvEIdJBKj0ip2qyeDbsJmLI+fHjIu5aMT1+p36CKOET7R3vviJfGzyF8KGlzt3n4T
hWCdPcG64aSM5I43CbZSHwW2hewyGJw8nljhHRWCMpFxMtfQkwHYEZAPRYkuzrrd7zCTCxfi6NI3
Y4VWei0UO/dizeg1lFjrJ6M/QwIIZ2Ryl2xZG2V6vqy1D6ua9seyalEFNe/Ndt1mT5vA9Xyiknxs
8yEnLhUFOp/iKaRK8FJQ4dIJQlqMyfD4EkAyrXuHnoKNIoiLYU2PYyAFwVUcZcsOKntx9LXSmX2/
uDJgb5QfJQvhpcY6vc/78l9Ll15h/Wgg2K1nnnATzKTccQK7DpQ8l0qBZ7mN4btV7D8ASCVvnR0B
XHSWUC1NtYFxU6K45oXyfiLwKnRf6PLjDWAjEvfKx9XfWScLFDXZPslTmUkDHFKHb/CV21VPozY9
EOtM1Bz6nXejm3jgVpi6PoKmAsvayNw2KmVghY0Pgyqd792cgu8wtYfpfpNJz8LNOYO/Y2EVu1KM
WRPg2VLfQzIjvh860UXNqO9eM+vGERlofqxwJY1LPST2XCXtzQBjv57scRSgcR7mhJFnhDCKm38U
qBRFLltXaO0BkrXt2jypFSZjVuKzBUwZ/4D4E1KkabiYtPD3uubPX8ZWi//93S8faFe5C1L8f7Mh
mYW2QU4tL7rXZbokbPmtqEBMCM1tsn0Jsl8a65zO4Qz20O4CGLTHenqp9oouT3ypvFK9bS50+hTw
e+e6O2dDdVcbrzLCl37d+eqvBqOqzhYMiWryUjLaLEgiqooazMOrduoedF+iPbnSdU1HYsGAY7DI
vJZlw8P5QGlwhW3KO7CckZAoRLOf81kspEvlmunNelayHs/aES1iWq2jUkkWl3NGSIAHtMkJr5SB
Yb6qYnjtfN6cSzIZkhMiqfWeVoQluFNIdqNi/jdQ+MZ9iadwSr5WKMtq0EnbTNbzQwo7qVUMKH/n
fqf1HI4+8jS1ZnzTr+Pj4xtDqVBmHX9SfIMhW1AMuYWC+KJJN7TNrLaHUcmJpskkuhp1o9RxCFqS
McNQIPfcQzANEmHocNH8xABr4Qs90k+KSPJGhqigdzIW9Lhsa0ShvUH8iWh6NXpreAPq3x8vFt5J
7VdeEvVBq+91k6KlOJZQk2SeARm/V9E6rcFfrlHkSbPq5QCootAhLDUEBogwvhCHnAKtxTxAHVej
kpLVgKP9+IeCLb23kwRv1xeiRVUPGHfR/NpLrUyHmTq8KCpE74+U2eNlkgyWpqVpKVztwOpFXTBu
qnkRd4blW4lbYN42dJ2blo4jp50YWfPuQqrc7DZcQfnFtyGiV2BtNTnUryY/P8zonQbhsLM1TShS
A/uw2Hgz+F83XoXnQRRWhbganE0fveGgagvcg3Yvt8C1hrf4rGpXqQk5EwGmYKy00b3W3kAzo+B6
9OLbycna5l1A0rqLvDC3fFHAY3BBSDF8xpM7UefT0wF7igl2DDwoBZnQotE0WZYTXjPqrbUQX3Sn
SG4uXG6I0Dobn+uitEBp1w+gSCJSr61nuPocLeC2UDGsdhBKZhZ6QCal6I/P7dmaCiDnFvCGkS67
JDt8WTKzmqg3heSe4ldek2NXy/yxE1MUhwXxpttajG90mNc/9e98y0Lc1iMorPTcgIQxM+28mXIF
n+rW3BNJZj4A/SCo6m2g9pC4HkfhTJ+MQiDahXz6EOFT9KN7WiTcDPjGEBjfQrPpfIJrunXd41/i
YJO27m/yxr1drMtWmcbt3NhakEBaz/aTEEXoLMFPZ815L1kGJmNSJqr8JY5ufaxWtRABV9hJgpNt
K3Uv24VV+WX1MuzN3Qzz3j2Wi1W4hluN1xHKrlek7YSlQ9DQrPfzpCqj1zzm3Zej+GhAxn+JFXuf
InDOzSlZKhLH6ZIW8wmla5iL4d1nFWCYXrJ8TxYTq2g6eeYEAQWHGv3e7lz0UkeJWiRvH5yiibHB
kx0H8Ny/XAZNWJ+qgrLn3Y/3I05MrxSv8BZmQSca0ld3vkH10ufU8YqLtBR9T872ojLhkPZFLCEr
ORgGTWlGBmHXBiA10STHkAgn/HqMhcJNb8JAsIWpLgvS4B/TEngV0B9SVmfjbBzanwNIGbBLNaqc
yS4q2oewp1kw50QzXeOMBV2VW+1+x/id2Ew0Ni83tL5p3Vou0JxtYDpDZQFT1JKvbkEL47pKEtgk
ohge3IPcnBtRaSWHz8XMc6yGvGeB50X9GKzDGkG0MqQETdvWRVRSNk6AfeOreaRu5FGKTT8an7cD
BG7YnxMW3OKCr21oeGndyzoWpBb/sm4mVMD6hOalUZhZOh6x3bhF5L2IbCuIgHJGezS7bkpaPGOr
NseFRpHn7OejdH7QRSfhzucA+94kvP+5B/UScguWkQrHNoaqEYWGNVZt4/AQdQ4PCWWt1Jy0TWRO
xRvWFx1QNvSgLofES1KSKkLBXlJo6c86wWVPMAiLJ6sfTWyBtvZgi247DKI6qnfM1HeQrl3MoJmP
RhSiNOy1zBHx/j8hcsR1YHJ+0C+2kPZqfUtMzPSaMAuYZBdNap/lkmKn4haG47+kEt9bLkDiqjoN
2fD8X2i8IeHP4pCAWs4abxYNHutCYIKEzAg/dZOg2ItM1PiiyPqNPC9jPJJmno0O3an9nlQUlfoF
0RkhS1MJFIjxsISLNVhFYD8LPCttPJ9ERRSVS9My/FsfAFNdo6PJOnsO04tJDne68b7xZf4qha8Z
WHC7XwIrDTLMBmZVAoVAe1xJzGvxAAO+yxCXBK8kYOgKt9PxDuKwgh8XsMmkFRTQIMZr623PDztL
1MqiEACtnvn8gMVCwI+7e9X05yyCReE3VMrk3a5tilSJNBkd58Pe+Q1gcHL+Xsb31oaj/mR+Z3k2
LuPiYuIGDCmDDsTJeomN8VTZ1MZbv2jNDjqkrR1KDxnKtfq21WncZyMZijj3g3f/XUAqWM5rw3lL
b9PGgtOoZ3BH9XQaaJfBY8UjutWTXXoUroyd7lwVnQWL7UJYCSo4f4RQTcnyS7zBg3qPa8yCoUq2
wlk5w5n3hIair7obIrRtu1cYZJokXoMP50QuKYo6NTLg/aw91/c/IJFVCwNor/ErTi92OVzD/vyD
k8b/fgPq7dfsqVHC1aDu5jBUhUum5vOHRCv/rZcP8M100uAL9yRhLDVr92qGTFSTYYdHkAXcSp/w
eP6FqFLrKJ0lxP2PDHtUwlfVCi+PR/w21BGEd/wlf1CMH85jPXRdS/g9uf3lvl7PMkwxeUW+ylXk
j8ggkGmbawe8jzR2gryRt7QWCVKAAcADbL8mtzkFbwD+d1Yx44O7mOvuDZI8bPp7G2FiRCZD0akK
+L0E4TiEUDipylGWmpXimExmmmFHIo4gdO3IwkeBPQtaC/eALEifsyxIkzBbpClaEyYdm6uMaY0u
nBsQqYhUgnOzlZiU+R+8T2toJ46UZiJw7w2BxzD3WkhYxjO9K+ndRYSTNFEaTPXMnNVqszPHsBuF
MU8nPfb31jsCYAtBoT2Dg+ZvGxP+3xqYJupcufz/eHWcSfMlCFgmQSXZz0tECeI4F5Qt4YZi9ypj
iCMjAbn/vUG1xv6lkh4QBeUaAb3/LpVFRmycUzalyhvKiZ2dayge0q2UvbnPp/wVZJPzpz55nqVA
8Ugqd+H5dvYggwjuj1U5Nsi9So5nobiFEFnIp1dUmEqaO0JaAPCwEfv2p9dPnHrpWNCRDeqKK9eb
+O73sSzZMCMhKrt2KkLtwb3NWz3N+341Rnbmvs+kpouPm+yO+WsEp7vSTGU+sRJePV/3U+enuxNi
wcW1sBzUKVVSrahw4aqDMTveaIFw/hGeQ0L6PPqHN8c9FZryDlVNbLSx0fI7fojWgjH0iErts1po
QyBV6n9NnmWhPdUM+N5z4Th6RlQXwvfdLXzsSdLw0jTJe+M41weAAUoTG89ZV7XLUDQ/SYQuTDjf
rFY28Jkrr3yidTFK7+wnW68gjL/svBrfAHdgIIKLov2rv6EN1OMnSdW5pqIhAiWHjHoLpH0pmpf1
TyAq6T1Kv5qjcVtTN2QIk1wAfDx+EMxCKE0756Bp43XJ/FfmM3/sWDIwMKsKExsbcuZ7H5m/KnR4
pfE7uIIEsSNkHAk22FKwsE3/mJEWKNx1f6Y/4QfoXLXJUXiz1X/X0K19QhdK7EIkGDJG1cMEchJZ
7GaLGEEDpflAsriM/EQRo0nkRP4ZuHR2a2Q8iGDX8MSposGa1LOI/8MJcJZRDZY156O57Nsf0SZ2
j5XCK8nlzWMCKBknGDnFgkKvdOHt9xF8Q//oT6whl4ntveH9JHObFJKYp565HHteKbbm4msMgQfK
P2ovhWEhV80E1UUdmUk6bf8FKsYDK+Wc1HtjTiQiwS/kOanGBRgDv6KBAoh9UIZPGcplAzYKD4jH
UVZedg8kFZbWiIiNkvDcvnCcQ/ZkBJt6adVznhes0C0dgVl/Bf0sH/7HbwEwdyvkp2FDv94WzgrY
HOPb0gkNvYSBs3S1/Q/x6aw9ctgzyIuz5JpGW5HlKY/sKBYvGxVKgCIkc2EsbGoIVzKA1nXOK+Aj
rl3o8KoXduaFvzfrDf3X9/WvE3hRK9egc6wSNDE7KzpB/OE179UzwdDgrLWwhhyh9fhrOWLwtjWN
MEGSXK64MGEWEO2L+GLrBGHDkDo82xWdRPrn7io+iYliU6oJslGKL986lMSVK5SGWwAFoulK9dg3
3neIwWkh64L7cSPdijVi8UHG7w41xhklTuU6ifKHqRuwDVHYDnvChx7DtYwVDiaiyKJ1MXMLDkS9
nAi8mmBqwRi7s7Q3hQAzycZuAHCt7YbtbK8STYgQvIoHlcXMR37q19X3dOFOAW4k6cKGjVyy6crj
y19Kwoqk/CkRRRM5iBRhfQ7NXiDeaUIAH0oxB5QLGApiXoe/WjcdlfMGQfUqnOXmTjfbzWYLM7Wt
dx/IBKalGhwYtkL48INKh9+IpG5jLQr39zruoCGxCtPsghB/fHR7USFgYhpaQRSITK4jpvBk7Kxl
PQOTHngyvsmK2x0cMnPCg12vylvUrn5uGst5023C5qar0BqVSCzpuhJKQ38VDxsjh8qkjLBLySue
feirrs5t4d9YqO/6whO1RuvfpUF9zOgL6Rmt582oD/w5sfXeidhxp5bm7rd2Rn81S3cqnAsTU4ra
xx5ORwvHFyECJenPy4fYt0fs1GFR1wrTHDH31isgQPfJTpzJMBWcxrARPmI9J/Je70EnW/vrxDGJ
SXUCNzKiYTw23acJXhpAgh5uYz6VH7cEqt6PHTWg5R4qZjb+LJqzECS+h2DqrAx0lVrh9fcekR8M
09th2qcfhOQi6rEiV4AqHNHD+mkDpA7PIeJqAhd853nMiqLBSZQs5GEp/3F95zymQa3JDLmFhprB
Fc5S81hTbKvp/f5+j3SWQKH83pJh5kNed7lscsXFO2ChR36mrjYCW668Dwy4I8xdNbFAxvxuIZu5
293fQj7hAzNARhjjd5vpIyP1zQ0xUFO59BJcyXdBR6CR6560JZNBHXdtTipdo2n+o9Rvsc1Njrc/
E5xUA1T2KKYE1qix6Re0aj83v/q65hGsOuAhZ8D6YljUYTYa3LfN7tqmW4dMEOt6N+1z/FYOJoeT
8Tj3snSFxsd4OCYIpngCeV2Gy/Ej8B7cy01OeXTXucDP4MWMYLlKHSNaeCPbJFGGW0iqjCET1ykE
ya1+/0iLc7NEZY1HeYa4LPW0URttmRzXX3KjiOew6/GghrS7IuKjV7gZXGuSLe3iz2fGrxwd8NP8
IzerKSJUkG1sjfNxB5APzun5imA2auiI6wBZs4OhUbOismRzDzeSgmJ/uxisuTiKQEvh7LiyPblk
FekBX0ySiqWqcAtIBEf9ONJ2DFCUV4b7VBWqlxKCjM9WHafZ8Mwh2pvca0Ugemo4CcPXXzqiFLN/
l0FtuorNF6JwpyvsN0L3RaUGSGpE69uGfMI2QojS1cJbPx9CWAkTkQIx6a+YhBbdm0nkr9S7Njkj
7ASpoCxUburL1isBlSn9ZE4MtaM7DD6ev4jtlTcI8R19VcKgZzrbp0zj2C0EajZ2FY+Q5HGhz6uv
4rOa03nOgQpwvEzdwjkcMkVwlvxsPxyqv2L5/SdYPY/KBlMbceZr/oG0jCTaTkqe6ioo9ynDhrlB
5M3A3+DT/imgrpB03Wh/WV3wO8FtbfjhbXq6SFNtbsB9fcaZXIdBcYg1R5umLeueG+firMTyGMo1
JMmdicC/i7GCFOFPSMqkUNp/Wt6sw8v0Jly//UmdBWH1qiYpMuvV4rPRuopdAEc6GRKbn+4WS3Z8
TVy3wN2lSNMv1/300Xh4LTyQeRoDES/rDJQ8Ba3TemFCF097vlbqfV4kjI/GfrfPOgrS76otJHKl
cZSdeDff1QBwHIvVzD66XERgdTPIoK5+wnR9FnJX4CaS0t1L7TZT35A6lxayCNAAjCgvo57kJZ1M
D4dWDHP8d8vjimnmFTfOedHAQ9VgjfPfomvlYByVOO2tGnGZ9TeDL1DMQnvrK6DhKe8A3Ff0SuDC
7lR/POw/AQ6e/NjNS5vnfTUsuD8DVFB2qa91S5xvUTO3pvqQrKothLpeZXo5l/v3qUpP4Svbx3NQ
BZ2yu8BTI5UTOQ+4vNwerLZQcbw7pw+27LuY6hMatg5BUFSxS+mU/+MUrbTyGfIt2YjI9dlJy7jK
v6v+D1c1GtiLAFnjTw0kwrYqLNaIaYwcYaYynkMhUMLFeEGpZNIUdSOkmUGSeL1kqhfysmRBTX1A
b8HS/Ra8REWTa7p2031/Zk3Q+ME8ca5PCsI8pFZpJs51tnH90Yc8t5XzdM5SpE+VM/VTMy3l1RW7
AwFlsKD3OXiIwtYXcbbbov96olXQ7frH0+kAdtKdCnfa4HonQ0zlOVHPaLyZ0JHHB/uHB4Ss8aSb
dzYVpotuo1X5C6HHCl5RsionQy1LHKUbZdPfx7s/bXjk5OqSs/K7UFz1e/Hzm6xU9mLJh50oX6YY
aE9AF8aLWF5YaXx/pwVqJ3p2cVNLeSPp3S6/NUAGONwcKgLxnqtnnwpwcNh8/UKqSMaOklQnc+nP
wizL0ibRrxOlBrCLcP0uBZ0CB5pO0zHyNhqCbkPwHOSQhnfMr99SBqdLeb/91PIK2WPtNFTWzjfn
0Hh2x4dZoJYo+3JGdjadYs2TNa/sTT+ptXs1Ev4wiYFd/S+SNeh9cfhVHc1oT/H7wWhvOznRYv9a
UVRpwnDtaXKU9DYekU1nAwiTOaiWFpU+ZfRG0s4NN2XrnUv9vdwHi1pbJwb96l0v7ONBN2GoNERY
FX9b947gpu9JEa0O0Tr31x8h0WsWd9Hbm3Z2os8qlUg7ciqBHg1bECnDarGWFGF4ryMOgfSoPX8f
IHgcvPpv8fv8f471+L9FlEWSmIw1MQYYXB6ziqhTYuLYCz1NTsOrTJjmy0exSf2nmKSNIIwUxUbc
TkeEbIDNohGg4t/QUBOx9IHwWNnCiy00wWf4NQbQrOFZWaYXvPY4Cpp5/a6p3ISDeiJ1q2ty5dBB
VWLPc9+56I1xU277m3mw40vL7VLTYk7gIyTjrObapmQcxzJqeQKAyFEGwRlA1NXm0/qUfP33vbF9
+5AcBHVw6MVg9DAUOg/1vmyJadPn11eiLSmkdaBxgrEVel1Zdy4SmviK5Y1VXMROuqvTQhS5ZYBe
sscwzTDKVz2h6UpTai/qzuiv+8fr73/+dj3pLjzjJyMqHMgnL3qcfrCuOxb0x8dWpNG5N5055iGE
s/e6PwNIJcHbyK58hMXNuEx+aZKWRNYenEv+BB3WksVxh1aj274D0Pl4y1Mhi0ICMrigqcguUwA6
dU7ZHEZ2PPJAytblNerC7hft1xn9txpwyQJ80zND5UXZBqyvojlZbTAGcHWRlls6d2PcvdfkiKHH
+n5Q/2xEOnlKQALFoxifZvRVnk23FBRGWPfvPSguJOBJ7fGfvI/xQ/1XhshNnkbHfo6S8MU0AC35
RMB5AWSqIbcVR1zoGZ5Lrp8qwcVLmKLr5e+NxoVRrqLrF5u6GDPSSA86nzjJgFf22tO4nSZ2YQsa
J+xcKyhIDzBnu9wPEaPSURTtArLQrJWajo9j0TnF6rTCj5S27vxIVoJXiGg1dUWN6p/fQbOfsgUj
msCoMGgTdd5YoIgIjtNeaENbpMQscn/REkcKkp9qdRkS4+VKFhtFXB5MO3/PXNoMjFeypVm6UfIs
QpEOw8Lsu/KM0qK8H7suas2gqpp12oN/2bJr28Ec7InLG62VbyHVNSI+SQ66CQguX/IQDhUvG9uN
QAhA7q9vGfKLJQUbFWucM6qXKjpsZD7L4sPOWYkCR/e4AunoZwlKhERqH6AR1mmzBFQo2NQ8ilqC
Sg2swj8cgQI/SbT5x+Z3pe2KCSYzuRyOkkRfzQa4/1k/NdbNUBG3fg9I+2WErECxKTaeyGxL/iNP
8exJ+MQO78GH0dKX11Fkc9oARNKAXapigaaQIqHowTZAKytKvv2LffysBlVLgLUnSoEb3GGWg73h
sded4DioExh6ttFT9c8+TEN2a5wrScfOM7sNS8amsv/q+YzbNMMJWEJ4oPGH6JkHFz9wIqFL51rT
2i3hlTage84vbwv+8NDesaitm3fW/9mQDvNrpg8TpK/bhu4IMng1eVA2u11KxZbgdlJ9iKmw7ixC
IjufmLbu/ayvvV09RL6wi0tUfeizXm86yxdUoOtj5p2ckcpUGKIJ8/vjSgkfI++BsN2dkIXJVH6g
cL6juIRyc9TD3D2FW8vRrsFIRi2bfRCQEkbEzvb9XviF0CV6BI/H2+9yxJmAswYUutEBfdV3EPzp
YPCAoQTVc0zdKvs0enTp+gWC7m8Z7B63rhr99ZTstN2dc9R+0iG/LaV0p8Qu9d9Rq41vyg4duUdh
wS3YGvEN3zaTSslzyD1Dsa0OH7PRTwWaHHDvdpvI4T2yi1+IjVjwkIpcWQBiXMHxp+Edcdb7Ial4
BkBivz98kZr7iDD3xohSKBYiJyMDyGNuDvSveS64wMCFGWZgXTLYmCtyo50OWTnVXmaWe/dDTOMD
TB7EAZ8I5nDUaDyXctNgNA2YgfDmISQupySaLr+Pdxk+9ztUx2yOIqz7NhsHfpsE326j/omZK68s
puXGg7bxVD0zQSqnyV7QJT+smbqgLoMAFX5RY222XZP0gtIOmfVx5TREuBdd6BT7f4h77ULtOpvO
GoBtlD8kvMoidoukuL8bAMOAhEcB5IhLRTxmm8g2FpjDqX7K3CdJeKQ1DTZppguE42RAUXi8xgZ7
9eKdjp57+FPv6oU//n0pB5ewfKsRsRoxBYFirZsAIEiG9nVVarvQ/xaRY70UQONb1Szrt2oqj4KR
g7QD2Tj6dLYlhtsYyige+WDGvy4Nsxjw9t2Q2Hs59YkO7ApE0RSr+j01DqKRhMLxKCW6cUcb5ng7
xUoRG6rtV2UYrwWXWKhYmBrvZj79u7TTEVSg5P9QL0QfsvttDm9AHRJM15fSm2IXIl4J2ihxROHa
TsJd1jdugjsGTJw6hjA/E0qYT1uD1cYQj7YcP3pAR3UR8Fvr0M4yu0Ps7yX4sWBQ+gt96nXUFLPT
NcaxIG+zku6l8jM/bRDIHIDoNbuqQOk2iS+U4QErjT//OVDEvHtve3umGduSDfQzbZk55FQmdsa2
i/m3E42FRxnHTtMgaxwncA766C1vMxl5+WJkR89w6XirJFfkKry3ShX0z4fL6PTgYZ5pEtgfylHn
p8YKIkWtykJm03yLdyTbKuBLmhXqQqSre/btHEAf9tFzNmj3mE3qEqTYN1K42/OeZOjElkjrYlH5
+6T3SGZOoq0etq9/pw5HaHQ76IrreFbZDk2mMnfrolJMwL1HSsjgVb6/sLIwAFMy1a+0yyol7eQo
/3lqSQvyy3Exf5rP4/bWmE/1C2mRKnQswLOt4QAk1gxLMrGjUt3Jwk1ExEiVjjls6INlboMPEreF
bcZ9y0cg09nHFoee/hlWinBHuJEw0CdXG1ECdNVdNmHVP1V1gywPJiUWaxNTPOErpWhJ8BTEh43c
rnN0/vEkhb/F/94RByEoE9fddhpRYmIZtP/ZXhL/PBZCpWaLADJL27JsG8nQrcQRJzGCKW644PP3
jDyC2S1yJt7hQmm2Dkb4tUsrpbeIRXVOCrmcJJ6eGkGF/ZR5rD679CQruYy3dRbVOAnyqpKojncY
SKy58NSpxsIhpW+D2PPyDwi0M1wjp/xI8uEyMljA+zrgneCsI2Mm4ZYbh3m7BIYV+85g6Yg01a90
GvADd/oguv4ZkDmWAs0nX7/5USm/xYf9tBtAYt/Zto2sDW5iVZcsswqTn0mBrzS89fwQ3INRXvDJ
U4CJ7IIRzxXTfXiNobJzFnmrYFt3lVt2bBI1KEwnyfzQVPYMWpjq+bo28QdffHgbWapnW2oOLu4+
GCjWhLkhEM8siB2W/+jq2GEaJL3OuLZ01pHP4kavkRbjuwLalRmr+QXE4jpLPoi3H5XAt6ZUCtm+
zQ7FYmfBbdQHAGKRKL3aBIPUtobFCsTvrTiH2vBwma16SIrpQkbQETixj7AQbgoDNEjQuiq6Y/Sb
ApSKBe1Ss/qRFLU0LsqR3aVihXCn6ZmelkfqmINIGplDdkJxgyNaZw0rq/Uo51qXgTb/NeumSuM3
kCU0vdwLDhcEAYQOzxf3mkZ3Ej7vf7tNg6bWKQQW/RjU6lJWPRmTng0ddCmKduSzm8Pcesvx/3XX
XZgNf+xWmmKrkQHn4JFczFawf9A+wIRKxZdmityX3rQENNEI3gM38mzAqQPbQ6eF4+SpBU0Pr7WV
D1xUAiqg2E5PuOv4GO8S1WtTf88eUWn4WevJf6JooPOc5sWh1nKVNsym7sQiCFpZVjQx2TngI8XY
2zgeo0nwEpO90P7NhtNTHSAO8gXEbasr+znSgGs+TQWzajQUaA8bCKxIN4MmdkO0xnzzvM3STeXi
Q/1PJQLOF8keuMagzPKOWKoH/Ff2MXkD+081LEb8sjxFlkUbccorZua35hPpMQAxtvElYY3vEftK
g3i0fREruf4cEmpEZS2KK+SNERtS9P7xe8Lx/4efVnmtd9Jfz6xH01j0hRxYsV0zMNu+QzxqN2cO
zirK4aTCuv45QEUOZFf02xwp8q7sWd4zy/9RUxishZmSqsIU3TrMD3Q5Qmhvz2vITXYrydlaWGke
m+IpBcsO+dvusxpKEL3Q3ceC/lK1q/lvboD0X6kSKSRIljVzRCV5Z0J9qW5Sv+em+AUxxvZCmc+Q
UqW3hQHleTrE32V9CkV3a31pqxlmzHwxew+6jqSbWVrEuGRORchCX5EnwC1Waxn1ora+SS7ooIq7
+7/hW2Nk3YPMYH8XL094d7zjGA2JAOHiJPfxFUvPgJdq+EdMbQeDTOXf5aNtn/E4xA28J482rHAq
GE9c4YNSo+3zX6stw8oJZGp88Ivg7Qt/pRz8TQt+eKmEkaBXR4/4EMqMzinJZq2jVjpttnghjj6K
EvV9dbgOdHhlSF3hYAGakfJDyxUB9fYWfan4xST621NDa3290+v/iJczvm2ErAik8dg0hkkxt1Gf
hcs2dSQnnUz2FlDzeBDgmrOcCa/lAIlpmryGCHgY9Cd5Jq1P0SHLHngJ+xW7JgVMqDuNGoRfHX5Y
yHXKFahp/sSlBVlQvi6XXbUY1McHEjaFH5wHdzZ01JFC/rJphNdh4hPrnwqwx99hB4DA8OvQ631o
vkAaGmRSdt/i7dhyilT8Wv3DeR0Ao9VdblahE7N6Erx/JdfQMbY0mWToxyMYdh7I1YcE18T7Q7WI
QTE4471GlSzmjIwPeysfqOZkSXRHOkwflRSU6LzjnQkh6N+Y+wZ4GBhQrUqw+fh1GypDmJQF7ANR
7ZemAQJSfM5pg3jJaTI+mhaQxJUKcWi9+F4AcJej8JdjZ0hGMhJ6K5te7SfQoUWmfX4Tf6CXKZ+s
iPQjajtse9XA8RdebYtwP5q+azNa8/GWb7jrkve9oKduAGuWGQhJAEFD0KWmkK/rrdOy4hXbiwvH
OIx7dIsuZDWOhd+5gL1oSIWJolwtz2L+dUFe3yosHYJzfO4j3gnikcE5tjqV0dIFWLpJnWZcvVxe
SHUSmNeXJoM1wKMFO/+JU7OC4FItZOZ9Z0zB7LuzqYtrA7OHIskKxvlSfLyOuRFzZxdpCrb/YSiC
9uiz4niQN0fgDARe9W6ylB24bX3/Qj0BI3OpgpRLJ1KRO8ZLGORVC7dVbJxs4lPTyPJa84JDhMoe
dy+C9VPjl0AInsIJa20vj3iG2KNBwDGNecI2Q4rihw7c44ehPrdgQpKU47ncHy5CzmMHXrOT1npp
7L2sTLiPFwg/czseoosyNLOtfgbqG7Q4gK578919cJXBm7eTtB11WMYy6xpSs/s0H5n4HCNH5mWh
iTb/b1RljRZf1nw1LjWExmWE7WJHZsHox0Ij0TYVAIBIPgk42ROWFHMayYwp9K+wWov9bRPT2Bqq
Sh9Va5pwk8OGOuYZm82vKY3EEmnI6AB6dTewbFLlJZfQ1IG9CQSMsjCN0JpRs/yBa0slag8Xv+Tv
hkNSSTS6klflLz6ERkD65zbb5qiaX+NJr2+og/W23n/TA9oRVtSIk2ujDRRjq8SSyf/QhMtqjl55
wKXeot/HQf9boyQ56lQYFJzEPOdiazuH4sy4d1flZsZaynG30G0EEosjeuI0dA/GDX/wx6mG7s/f
T4/yDNDksPB7m6e5maWjdkADKlDi+5FQie3LEffweL6o3j2qoMOEjy5H6cgvFdFpAq/nEiqE0v+a
t2+e5GDuqt46B2IOAgJLImX96RhVjh904JuwI42eCR+hRr3Ge+uB04rXN/ppdJzVv6nz1AYQDtiS
iw46LZjT10YZXZW1hgbJ6oLZLfl7l6GxSN88QeVrW1DvluGlhh5nTKKqY8fZLdoWhvLzaZ95FjMQ
sfXm+ayRI0E/XkAheHmavTB7LzGRSJhkEi0/H7UARk0vO795jRiqlcpZqHvO46uiSxdfMamKwjRq
lVzlVLNsqbj0yJ1z/Sd1OlOgS6+Eshi3p/pHDAZfvCVk6ikcG0zUwvPYlIhDgT2CtEl/j94WKCVi
iatabcULVyTUG3f6ebnAYXJ3IyqX8KAloypry7FhTYYLqPMfCrzllN11eR2CM+yUwS3cMMioZ08+
9T5s2P6L8Etc7mcc7Wlhz7K3XBWM6/zElgIOs1kfilpRWwBv4JPMD/ptSvRTK+MoVinVa6n1Ag78
ipYEdRH5JIq59uYovLHeBirXKQiUhoSsQ0oxtSM6+G9Qc9hBJFzw+yUPN5C2O9k7NXJJ8PaE7KJT
4k5dXcRLXdJRAmF+6LI7OUYRnqzs9lEkwsp+92Q3vABmeyoL/+HTJdoBoQ0Tn/kjOU7uXMgoL+Jn
xszxwhZH+JdTEHiJsiqCb1LvwHE792vwUg4A6sI9pSllAXa+iI7koZjxQfRwHIA9Bd8ka54jNWCW
+9z1vVJ8l2Us7cbaF7Y/ketLbLxbB3mFkzIzDbeo175lWek9UySM4xFX7wcLw+E0ARXxl9GcHfQt
T0pEdXQiwICuT4sxfldffdpJtIgZ6fRLRYnBvK5zustpLk+F5L4mRUSdFEw6C9GXaLLA2OyBQY6x
MIqDCT2SM8LTwcJI30bN83Ni2SCsdiKHzNbpwbrSBbTUPG70LnYI4uVx2G/bIpoptmy2cAWNzYku
IaxrszsU2MCyYESCVxHhM7XLOo3MaeaLu2qBvy/KNjQZ5XkYsIRDXglt/1+QHb8jzJAWn1Di1uEA
m+MQFnNlaRfQZnXx79a2i1huReT7NuRDzk8hgdNEiH+iysdWdQOyp5LdwQjayQEWHxqKLVYAS58I
JxcUf2yDsA8NNXug3oVMii0OFnvkxM5qWG3QiRrpI422GKhGG5vlVkKkykSawdpxgqgPofkxxyh2
2wU2kpeh8D2w9ivoraNJU7rEEVIdH1F585kTMhjseqZWyFHdETpOYes4+SI2h72ZWYHGvuBjX5Ke
2A69Eru/B+SVbeV4LyE4jMQ+8QrmnGNuU1Bdru9cKWCi8G7kO3FKVIkt1u58l9oWmfANql0KH6cI
p8hFwp/U04w5NmMhwtgmF8ztFgmbZXUtrroG7izsY7y6d0mjM9y+Z6FyhswXA3bSvMMSuiam4oaZ
kP1xuztDu9HGgj8A6KaKuBu6TR4To1dIM5Fa/0H7H5WBXphigRAyEzO6wbUzt54RKjWQbJvGr5Od
ZdVLLPeqDdPI0FMnvSxU0PcPE9tcr+466z/2aRvDmGsqMB8rUwrOKz/edGt8h5mPtqxVL9neu+J/
Rk6kKfAjSu9eWgbKmeAOiHfVXtTCd25os9k2CGSwytMmxdU6/kVQ9UO5lye/un1yH6n7UkKY/Nfd
oX6W4LbqPqz0XI1NSO8btTCy3d6ELoVtVaMAZk1ELu/X7AS6neYHg793xbEwK0MP85t7EfKY0Fou
/ZrWjnGE9jd1lvXVoxJ8DUYllReJBmyA9XULAD5ki1nFynmMiGaw/pqr9h5XOtXMo6q8FUpfoWUS
RxyIRGNY+XtEx00uVMeJVIeB095OF7v41P7kPY5BlSWyDDAA3J3nQbliJV4iGxLU6JAoShF0Coeb
WydRgM5i6JjjAsXYM6JXuHaq7VGhGNyQHRhMpFCLN+iF66GERkVDhtnDonGqpSEoXLN7vQizVbSE
QeiUIeBM3hwZ1mJHRtAop9MdzUorGqAd7cBqJyVhTNjiDiZwq0hsU82066geU1/OQNnISaunPysO
lbR4Zv5+UQxgCkcaHOZnTo7keo5sUWmbWv410S4RaWAwyAkAZP8jRyA0hyQSyNT/k+qr/UM6Y6Mw
eHbzFOB+UkuME4gXAhjGpwp0+ju1AlDzIQVqpz9QYJ9IRYDbUx3wOFQ49m9U5Zd7oZg5aAUrib9x
zOZot+Gw2nWF75fqQ/Uvnl1s4/12GhNBIauwfyETzujBXxkDguZE2uHzeuo1PjxL3WJVFF/NzNdh
4MLAkVTlwQanKtBVWl1i2XXRNOxWJMoy82PDnHkLRojYH8uyPi/AurdD64+C2fy6YxO7PH/ZB892
Zm/C4Kqi0ojmHi87FTeYFfWQSwpH6kpInwbsvYedwAbrdmeLCHDV5G4UWJXLxLI6a51xKYLJJmpT
6dD0DR6I0i/ZtnIwOuxz+gaHWLHwQedXE6o0BZlyrIcA6UTHg54Utm+cnfDt3uwZSxU27G74BW6z
rAjJCGTAaZKlBb0nkhkcoBlvJ87WC4fdvVdYzz+e1UHhOBtbKy/E6HNpqMonKL5Os7CvpBgRDC9J
AfpQhXFcxCZDtK/SrJEuDY4c/RkPKzg/H3qHs0qTE6lYAPxN/aENjuqbbCamMUsKEwympyZn6dSo
HAYC1chBvimtzduCc3c/C8BoyMMrgS/lMZT/2aJEzDqnbKJfvygx1Y0vIVYv+ZksXnXOT7+pkKGU
JRZFjLlL3y+SVvwQ75KiUj9vXftl3+AKr4uYSg/rifhIQmYcz/JyooSp/V8h2yR129PT15CmExRQ
XFCU75wCi9nBh0iQZ+MC/RmjyIPsqZ5NzcgkArAMxrap1iC84tFKrjN1cnElXBHVBVn0y9DO1RX0
MMPPzyO2RKGJm4ibXUsWciWXUzHtD9DIPTIO2Uy1W3RPI+YKvsCRuC5j0AtueSgm7vvAy4ZNCXjw
alsJTng5i6bJ86cBWXhhd2xJ65gak+bp2jbb6YJsUh7QVdwYBur4lRxhm31U9AMB4Shxx0A1aPBM
RfZTqrM6KLNJ4AedOMEdd+c9pKqvM9/Thv2FXQtSshk1g+VkPVpNeMsFKmzZ0mDdacOo1sO4MaNA
oCjbfEi1/+G4AIgapHOJEFyTIImoPVoz+7TSm/HJPO4KO0hTWVAbSrg/uJI7HmcrIRks+pSU76Wj
r2qOHzEfF5EUxpNW3JsDGcx4CZ/4swMSPH0pnrO+DJwJ09GdZLNhoh7DX11lDtgGM7xYlyCGeJaR
/uzDCKsku4oLYASd8fppW3+dYnLEn4ZEP7jRoOW+mUbLKrVLBKE03ox/aZ7Iqu7u29miOpNs5pd6
xxohwB0+kL4MQaiI5hEk3+nj/LwfqzNo9KrT6SO6RQVNGtKenEjZQz2GyxpUfjrKFn/qKWHm590A
lF8eW2UP8Fnz57l6+G7Mc92XfUliVeafUIYw832ZMNziafr/YVozKR/nRO5G7WgwMlu1O3h37+5r
KTevhqpmdQ7L9xAK5MZ+iCH0yVNWSBYUcQvUyogdtcI/XZUpmFwT+esdVIynxqzZleyl6WWm8dmc
u79eceM6H0CFDkSLmKIcqcqpQJ3Z3Dptqv4bDqCf7MAAOs94uC/6cHYzHJHK1zkY38RcUoFvrd+e
mYdHu1dN5ceCL7B2lK0QniZTXVDJR4edp8r6qHmg1uruBjze08wsp2Fap/csDLEI58pMjv3cU9kR
umL/DB0dwpLiRxmbdU3uCI+AXQ2ZWLnC+j0LGjFcb1fSbCFAHrj8m/Pbbkg3EfLOw3XRngLUM5zm
sQWfbWfTfaxtBQGrmkn5P9xzr9MlA52AyXAeJSgdU0+sSUlh6dTiCWQwGWVIm/qS8rmSvUHgT4Cs
8zRqmg7SfUB65LlIL10DTt12ccnc0DrRrsDU5BHAKm0sQgBNaBbsLbXxATxNjYwXfrVxGV12ZPiy
z9rD86llJcY88ReVkuGW+4vtmFkH8A3zAHU/fk6tgRsm4jJtRfKzwwUZZ8ZqzC9bu4QDlW0DLkY0
Pqbl+FoJ0FxeFn7srghuCv9WGjX0/bXtQ1m8tVN3wr+lIudGAjXz+t9rCHwsaQ7U5ere/Q8zFbse
vH80Kp/n2WNzHh6kbYNIzWdvFMCeLCxZBAcJ2HXAN28OhtpDbSbiVkIyWW0VmbHO2WgwjskjU4R+
B96A1RQQ838e2xAd3dHXAtkp2rEArosHI/mewpsrRvxW1WAWZFyHr6QqvFsKoO9T7dVCbyfEX91p
QekvYFlriVy2btM2n8i9xzVEYfRa8plQl492kY8l8U9jRpBEpHbOLwhaIQWtXM36+moLw4OGedMH
p6QXS7jObs0Sk/jVpv1lVGuiTCm1MyZK3McQtKbZK/7+4ArY6P6+qVg1BW8hezRN77dhVbgHEXX+
BhE9ahhDrQlNi3TykSIOnW0abfSui6wRWs/TU6tR1Dl98V94Nqhy9wO1mbsvXCunHpI6jlPa46my
5WiKyLYl+K5j2nnyJI1xfJCYJXNYLRLPtkgNxub0gCV50Hn5FlXbY3ZeidzTMjGo7G1h8xvyTTST
wN8UpR68Xl/rKtu44k427qriOkHVnrvnpPTuFO5ZagEQbHlEPjGiITy/TMi1gaqBoVMtmMSCAXY7
DWcwPJC9gNesZzTQvl9JaV7AC2GfWP/N7p9thQtxZpxbbjcjDI8Fohdp6w3tm6MbAWnKNCvAOrXU
Vz/pDc0v8W4yWjnLVSZh+AHsM/YbYqqqYokyieaTwZWz6U3RbIh6lubnFWW2Z2KwuNLiWIb3yvJy
5gQGiA6Rdi7AlKglniaWa8NEqO3dih65Z36XoCWBmUgca4j90JC9NCYMjRTvaZbaQQSjBoElC5K7
5NrEYaoJcVRsxqnj4/ABog0kg6oOh/8ywO29xkU9lJ3T+13GBjNM2enVq8lIkxh2QHgOhp2HET7q
THujUxUSkYxMXXQz7R2Rdi9WaGAnWwXSAiXoN6cJrokmsnan/YzU97R6PgiV57OlzHqgAoC6e5oy
npg7gwQki04zeZ3Ymj8BZM9cG7ZOWUojO/eshrx/oBTAeDLeSVMLC9w29675WhYE9FyGhw15avb3
q0pVwaSI1nEt+Uqc5ZqL0ssYSln1NkY2iOAWj0N24Y86FbKslFSG8pdJjWMyIlVdzLgQiVcVZqCi
QgRrebMSbsc3zzs8cQthqsLV0x7p425tS9UGYsA4Xzda9sA+3vRBtKM6W0m1dpectjXNN7EY8Pcf
Ocarpz9VCu05Ptku0rv8+0/UrLRjI8/89jtXIluJmKiE0lPfNeWSaS9VIykZhfCS8zbkJl/MRoxs
RwqZ+NG30jnLO8lUGn5A37RFy3rhVJMSwcYOUgty0zykPaTeJGn+cOIZ3qHVSpmWM3UTJNlKG0D6
6CGtH/nCcHyrqRu6JPTyg5PBKLW2PE4ULA9LBdX7ODw+RGfPtI99SUvOgXIeEzCHdDcmhqvge4f9
0lVWvLsH25yy1fcTZ45P9O0jO0St6eil5ixRJQM7u4mS/xEkuayeC/kcqWlvCu6OBgZRlqJbM7VX
oD5HEieO42OwKP8G1Oa0XRKbScEKL7WC4t6cLPVinvaVhWpsJd7BKeDI9EYzhTY3Z/lbakvilxmZ
3B5y75M+9pNZLzJnXhB1v+d25x5SJIdRRG9R2B15OlpiJRHmfybiHjsXtshmZqVO7U2tI1+Z7chW
BBMuTmNu4EEzvB/b5iYJ2rKuntXw4qUk3fUOdngdcuRRAbVT5icGyJJCKRT8olwwAXZpzfgL/o3g
Br4L6dowfWA8Fo3GfIU7PLdMeaG2/p74cGzHcAiwSAuCD2WBHaA1uQ2voZpmOdcdrZlPj/izNAMV
CKKw/mNKV+pXZn+zXU5ZgYncm+ajZkZ/KpSlnxVExU3UNTMN0wnsXrJ/BTXaGck9Ni/ZQU653/7D
Z3Wm5uBwwvDzfHdsIAEBDKbIHsJ4MlqV/bRunFv3bobIvAPnCSlnIxPVVs7voaE5rehPy63ukgrh
GXPk+0e8NfEo7G+y/UXlVpbj9aL2QWbLSvTHpvdl55Lv4/w7rFJV496CSDQmFGG97o7tRYTmOsYm
uCARff9hLMS6onGeUk9rjtHXHzyDMxcAa7hABDHyQsd8BRujBiKB+IEo7n6ChuhT7BkMNIUloG6J
y+ZtptzZ/qQiTESxC4xwnmy3VJJVf+ttNjfp/wqtPRVPt7v8JN/b+8bX8ybGr/NAu00ilUOXqewI
g8QTsDCxPZuRzXj/7nzuays/CRmJkg7ZFaeEnckecdSrkrojxoybSQbQvh5cFM/Ibazc/XLOlXet
KyeDo1GHe6+AqFcOtCvMeLVt5nkTdtKnXR0sumRMJHveR4AWE1PNEwwnsojS94irxgDZ0F6zeotX
Z+tMNhRPF0ZBVHhjYSNk/qSkgLqnkv4MPjyXoO3j/9NFDcVGz5iZ7de6r+n0DqpLh4IGzNm7/BNK
NEsesghEplzTIiub9F0wGdahTxQBiHnmVzlDYOQk1EhMrYauUPlQMuFys4sNS7g3/uiZI7FTLDgV
w0ZCYXoJYrttcetVr/0o299Finf8vTiDByaK9VwjDybjIEtTao32Oosd7WLAwI+nNokLT8kYq3oC
PF2v/SHw5CicPh0F3+XhuxtbStSOzv4sXb/MSSsBX+Wwt/3Zg8kmZVxw5DMBEz+uja/z4LWK664p
K6V1jvkrVGFTkvJxD1iEc8SEaba5vxTXI5OsaHIXVIPzA9YBDjzX3d4EtWD6WJLVqi9TrwkY/XvL
1OV5IMAXw8/XGGsBk/ijsCMzX4N5PsEomE2YGfVwP+tOC7TpsRpl1mEZYhBR+vtFfaMxvWkCUjRF
QvovEluJKNncYNbtcWElCd0CruLx/V4pLqT6Ii0n5m1BRRokR9GLIpYVFKxkz8mYeRwr6pDWTpFR
PiiFHLqzRNdHSu+viSbY87W4dLxqWo6/b+3BoIP1RO4xYSZioSQ94YNz811GRSeAckIRCXeoIiJd
msucizDnl++hdtvFMswFTTIJ3B1Sq8KY7NlMUUdgdWdB3Wxv70eJkadgHKeb2v2tTIi1fgilNvvV
rgBTuzOxl3LT4ljSR1FFGD/oDW2FRrcze0H97rDBBE4kMMLUqqQyfHBVaxBywvzSxtQpTf1n/+8v
ta3/DS2cbBbp3yp85ZEBFkgepJ3wl8CmNCkrngFegbzHf2JuT5tOxMk84EOyEzFml1YTp8ZHEJps
7rYm6VlQ8yS34KTxZhnO1jYr4Ao2xF5BLwZBtBOeoFf2jc540T+3FvzoUhTSjiZ52/1VheDVOPXI
WX8jdMXWPGf2HfcCCNtz4vX4bErYsad5MzZrR8zMJioCtt0gnSxvjmtt7L3NUjnOkjezBe7g0m05
BVjNQCAuAB4KV/O67xOzT8fDAtM79esdzfRK+tO7/CJNJ8IY5sSPKIWNzt5Txa2B3sWz72M9AXIr
DH0xKZeHVpCdalpH7dutNV44a47O/h6KP4mUzKga/tkGmIBy4Ui9PmkVYqq3Woc0Nuo3TpOW8Nww
8Tti93QesY/89XQqQn1z1Xe27d4bS3C7JyRyiRAAtyJYkqC9mw9uvYkIJnY78eS3fODQfGUInvxG
QUH+N7AadxC+8YvMvbkN0WIx2ReV8jdbYWM2nShn53VbheP52oNXnzzvw70KC6xJMQr6ikTipO/k
7ihGlqsT3tLmVuYHjN7JbgJF/eFO5q4PKSp8uD86qlPDw6bwQiQZh/0vFYbjyWcR911q1YsUGLAG
C6pflakhjGmV5fcd4byCaNpJ7jStL8A/UueBhUHAcAGCYIHIdLjiXaovWG3tP66ZE2xicS6hYqgj
1sOAx0LSbAUzt5rShDNnkbHmqwXkUq+pUY7aAoe+gIz0qfn9+Cy/YremHNrrxJtD+ES6GIlgtrFz
/GSKVY7XW+1KcGnHD98Ya5beB9yFHl5UJqh+29NUb0q0JxwGAuWGOWKComwUGsJjER7En1hViyIl
xqag6WP06SBGm+9XXdtzT+DCuFSR8msDjhfht+8FuDBx709vyIqwnxo/JjMWHEwwhCJApl3ySJEa
wbRwkqZ2n+RK3tEkNmt9zsUr1RMYWmyhlyrRK0S880NIW5DzkNi6HXSJL1ZtlQmCxadjbbvTMkKI
JybTd2fbyKKqdz+aD0kcXzXvG9nVnKxyv/pFcKYu8IgUrzSO4PrXz3LflP0A8Ona6Mt2QKpvzwXY
T1y52dLjkamTTgHF15Pj+fx7rtPfukFRFMZyDZ5M36ELYQG7jGFvGno6mzsPNs3EtuXkI0/76hWH
FyN9obsgNWpCrA/LFm/NP69cBIuB1DRBWS+mGxJLilCIxWV2tcK21R7jhuJnoLpcVnQ6ku4ocCI3
u8jHbkjGki8YYNmElPw7CZZNLwQeDR7DoXi3PAbqJQL7jE88Y84Da6H+NC2tZRSmI+M2c/PrTOdb
2re+GFOdoqJOWRJ5MhJTd8Im7xHup/SGBi8Dv2RY6643kh1LGMjv1k0E7A9v54h92oBWpwHncDM2
xuyGgJyhSt3S6urJkd4vYqme2s6LBt9Qxps6jGvNUW/V3b78FEkycDj9cenBCChBQjqHE2fSC9/0
2feQqm3KRXJ+NYsOO+I4ZLSuTQj0MbdF+H3WwuGoRC1rkEuat1wNDBwngiKAl8Y0/dT/c7QaktIW
C24ev0GnDXwbZ37u7VOFP5qe0f1V9xe+lLNz8RLnlVO6e7U9vlPxnOYfLuZq7wtzaEH7EozDZNI0
CFthtDBfvUuRqW65Fmx6dFFrAiQTK5i/aZayHa13WT9yaHzsTgUFzuRJod+/1ooEG3uGmowMu2mK
mm9ym46RU2a6Ck4JRf/OSxIr46gKloDXkFkd7kVb9g2APxQkF8zRpHOxAyvRoByxrT33Pc7KYflY
0n3rwRg3/1lULJIlBftYfhusIz835QujsT+ZAAPsGB7koe273iYYgJyZ2kJrv9WneQLGFxDPtnOp
AeQYvzYYwcmAvxFPPQ7GtVFGox5g6mlj0u2YpRREJd7P4AoKhbnGEITrYD6qCE4CUTPNNBnUwYM/
K3Vo3FV8csQgLgTps++1P7SHXrGlpM+x0uUMVoCNz1g/joJW8QosntKaCef+AKev1ZQ+Zy2IItw5
FeBjt/aRi4oYT6gSBXtHspjljIWKMXTH1MVTf+HrsJFV9hy1mMy2wj5NT5GDVJKGs6Hu7WVCHivA
fKkXs2YoShUGL9EdScVEusjVxiNWGylIGQJVN9S1jmMZchfApWIazjHrNt+dFalDxT+8OfLNAngT
HH6g9tuFATQpyQQjH4Rp3NVE9xu97IUbjB3uVRmWT8wTXcckebld4PXh0Ykx8jW+o7/QLJAOPafW
SIHRNTL0UExpVAqGP4PUJ/GI9ldJx4DznkN5yBotBkU7+RQHg7dnMB66rLYY+H18ETiR4ZZq8KEb
5yyNDyQ9+1jFbNe21bWjjLFd0bVnwMhmVMyCsx4gtHNeW5pRpvVGn8+y2pncxP9HdD4JDZ3wQC90
IiX44WldcPbrK/iwwrGBPH0fug4TrMOnTHg4TD8oSnrdHl2llC3NXdtF+LsEZ7IXM0PG2NvvOEhX
cvDIy/L0W0UZRrLXJD6AnZpjza6Y2HQgMZqHxpATx2TkXUUCPxJPFDHhvoYpZ38rTaYzE5sPIYrW
Q+Y1CCb/WbPNALl5QCOyVMaavmSrcGr4qKHHncOFv4I/kfU4SU/+SGilrJ3t9sb2+B2sSXWPhfLz
F5zHO9822RoBEXx9EYWAIBTGZoc9xfAbz4ENKyU2JVZSaKzjrnofS4zjLeZ4KvEZECUufL4G2UMf
4qMnT8FO0d2zUgxnrYdOtW1bB81ci6Y8pyUCjNvbqNfP6T2JrDw5mM4bSHZ5cVoyMP9PqqOZaaN6
igLtoMdtKxoFI+cuiorqiz/7cSZmJ76YDwoL1MxcE+9eE2Xz6T+43agTENOD8jd6de0d1yhNIZJW
jb0SBccHm32LCP1KPmZZdQGuz5fOfCM0H6aCsGodK/IrjmTGe6MZi9eEOyMgKUrlGVH3v2VyLOjc
Hf5K8OmuKzYgupK5s5IhvNaVWppYVvrTtfuo4tUaA3hfwcZS+HDUkLji+CU5cKdnPkX3mQRNDWN+
TYeq2DWrEOIm+F19Ip28w2Aimhghz5qSGNk7DYUdhhvJTh5zPoufhnKnDsygo0AiqA8qq71X+KxY
m0+L9xfADhGF0d+U7ccl2IGhMKRRtb+J3VOsYFuiiDXnqxOJ75TedVBhla4+Y+CoXODleGv8OfuV
pE6rnXc5AUgy+LdKKMPjDhnTn8qsR0yCuzKEBA/nSUZJyz+nMTuMXMQH1FxEAPi8xBBWWri0QRrS
tWabacz4Z6a2Mz5DhHC3JMopm3wUR11ufGKA1i7ER3/eNjLkxdYfZY4o0h3afYTdmYTxmDI/3yOi
yJyKEpgKgX/hyC0uMWi4ejPJGNOl7FYsSVKydQRqOT9BlaInMej6aBXN0VNHn1LzEbRQ+hi43QsA
e3FN8Wn/gcAmMGWksZUNdYOrsZISDykFtUejU2fLrW3q3QIe2rRgwcNgy/eernn9tYgyyaV8FWR7
07M2HjJvZnh3c/TLIj+lKl+9wu1go5nXLO/Kzp9TMxeqVDaR1E3UTn2kZvdUJe+NLPaTYopwiAdO
6nr5m4O1iFReps03Rhs/F1p1+bA+Ifn6ctqIeCdZ1P7zv0EphXlbCvGxHUeaYj7EnGyBWSn98s1U
pD6G8hwLZCjLLYe29m0gj7jnl95jLzF+Cey8DLuHCEXzQ6ZTPPas+MzQj+AQ+KUg3JPemrhcf9Rl
NupTGX9wwraRisMQTqSrvgp0YwcrDPDFrvLbLwdrbMOegRsruJZ6P5JzGKJpuuLZEKRizp+cZo33
tw4DRyJTGTcbwmjuREW1J4IhTXOySXsePIBVesDrQYkg0V8+ZlPJTTv5qncyG6RGgs04ibQh1csZ
Lz+SKEw4jEb7NFCy295P/qItEc9GaycFqom/OeneNoVv/XnMaz/x6H79FGnMxg8rSRj7BsCfo7Yx
s2wqthDroCw+tsnJgrZCc7+vs2S/8fP1IKRQB5oLDjZ3rF+96unoT6c4XOYeZqegYymNxNosto/W
LBlpvucEKcOQjCKOJlpDuegmTnzgfHR4rznlYlnFIoW+3280o9uF6PVCp0wFzKbmbICV69ZdFXah
ju1rWuyWUAyWKvPQBFNZ/8mtOIpYUO9UXMsuhNVVDCVLuqhio25E1/JpYfELlkwUXphVfqALc7Zh
eAB4g+Vc1yZAnJc6bgJCBglLnkJZpyE07DNNeHr0ib5zlMEHxS2Zl3NrferbM2unWkY77wVeCDqK
b2IfFQQMgX5+rwP+VoGL+TAWYLLPm0u36TXOnsJpZ7Gew/vv/ajg1JdfqNulBZJmX8WCT87Fz+2i
ed9Nh0UO2hSXXuiHafbVXbRYJsTl+uYfSzRJ25c9tl9qktRIfMy8RP5eOVRfvYdhmFEcPYaSwFv/
S8v43TSrFBrOiRM81AegZYXSy3dx+NWyijF9ByL8ZUHKp+4X72nwV4jLNNowxOFltZqskwIa5nbd
hSgxleYK46W3rvcpIJFQq+AEBM0Wu+GONLXT4SpTfERDuIoR1UV56S3ITdeb1hqTX/2L9LrcyXDa
pWc2DmmjrSn9n1mX6QbS5yQsaJbqCnXwMJIou69l5dF+ZJqXMH2ivMfAS6GQE27xgwEgE1PGAWu/
DMLhWjh+JAvR50t3lFuVpDWXJqoz63DDABmMzKKwbSJMr0CPMmt+q/1MU6PkV9s3kAL99D1fLPsr
KJAd99TI/JcS1+sDkoKEUzpDZyFwJi9FldHuNiUm0RBqngeetz4aIwP1Jw+18SUKouSFnp98iTZ0
91KZlXKUESxt7FhHR6KtAIoiH0hzf5VIeNxmXluvHCMFhut/oP4Qu8/xigVB+yxskiNZ+rlb/gYo
slvIUBTinKdwFBczqUrR1sGcGs7EJyFgw+GIJ5ol/VzTUHFzlCT3ATgAy32WMVeuVzkLSuA/8bsY
zcFplYNoyNfT//xkjtq2q/lp2cUa7a9UIp0Tk9VORMJTHvjCXJQ1S8ajUoaS2y1Onzp8+QoP/LlL
Y4pfVKW9xjDhenFuboepGMZuH0fhLv+QQlX5XyH6ZS3AKbe2q7871/4geIaCOcKWEpYMq0J0PUcN
ut88PXJ2Ain+XPfNnJyVO3xarQDftBZN99/Kr2bUjAd5pBiq5vHT+BBpt1cDw6zrYATBsHx1t/cq
zZcT4hGo4xKBkV1iviR6EYe67unYDroygUuKiaIcDJWC9YKe/8p68e2juzottLNq+iBcP6dUNRZW
yCJIrlCY11slZ/yfoHGHGpdwsgkNzxQyYGb0kz0HyKvVYC1uOEnk//wFH1tI5r5HhGPIjHe2QZ6j
ow3A2kpqltah5cd1Dxpzn2sLfiqjZvycZ5oNP8TLtYJq3jaYmx2n+7uxvi7uCNOb9QkdKr8UhqwR
n8+enV+NWprrBleZEDQ2MqsKbrqno67jG4gA0rJ75Lt1EZf8MXdDJXOdx+iMI158V1TUJRA9ADJ0
jexWoaPpSO7xdKKvNFhyw0p0KWkuSnYRMqa2muJWW/YBAaQpYHACELM8T6q8ODaJZTBlHZW0kkDU
jWnHD9icfV0YFyIMBllgTJrpxD9aou5BLVvkEMIQ5q2YloWUjyY/2VatHie30r1MwFztJa00OgNt
T8xtZmsi+m5rMn/UB7SGPeUbdrQfiqKe50XyyF32PZwGkc6vFRgv9O9BXxWbQySzzFA9XyPSBeo2
KRbFy+XTvDhzwMUdhKeH/4q8DCJ1bBtl+jWJnd/We6+o6FcijPnzoyLMs16gTUpFqcpPhRaCbqPh
PhJfZW71qw2+jhTPdWUTTjllputAe6i8Wla6+ID/Y37ZSdlyYUOQ55uHsZiYSVYoElMrdQdwhJNx
VaKLfCRZn6JKHW4/QC3OCOq+SlNROmBHlXwmsmmVfSlZj5OYtSArgLVgBGPlkzpmecB5OCKcZ+eP
eWJZFAOZujbc5mQL8DIoN5hmr4PYHVbNvtVqLIyv2+VL1t9IyQyaLUndWV7UVbCFMqfOgizE+PWM
7Oz1vpQhga9ndeB2+E4nmesgEwPnRMNVYsdfnIrsc360PFxmdgfYb54PtRKMjdQ+VIAMjtEt5Nwt
ujntqsMagkSXU1M1ndgc11xoQlrJnMv4cHvcRaYXb2078kNyLP66zZoAo/saVs1IW0DYq4CpQjSN
iRMc610g33ANOFmh3HyTp+PkMe+bB6wvW0ta9vSTqaydu0wvtjKsgQYZDb5sD9mixBO9gZy1LlMp
FAgKwxmqyDVw4XZvazcKMLUmFtpooCmsXqbEuYK06cdQ/jRR/s0rGI+kTc0b2zH3rDlU+Mhs48sI
KdA3BoIcJX2DPJ7kJVl5B56+xmZ1zEgo+taVs+xlc+OJgp2Sga3RTnr9hHz6RqqYkGDqHqpLS7KW
lrgfJ5zncuFoehkg3WNtYgoEzyXK8ejh2C41Z+g4BZiw9E/wVJnccIx+keeiXbrl0IZECSMxmhi3
GbOckoczSpAukgPx7kwOLgBHemRHqjTm87vl1HVz3rolQL3eNdwact6jUGFrARbmuoWsu6E5pWlF
iTlap2+DnGm+buGZsqp79v0xmxHdkizplxrllg4cSfvOR7GlO2h5+cM5n10JFTi7AvCoEo61ezum
HJDovR78fIRUPFAKJnPG63c0WlMUlgA/SUr+fe0wmCkC6xhdSCOeFNDWN97ldLRG1eELE+WpuCxL
ZvnUb+l8YUTxqL4Fd/M3PaYcW3bCOSfeTKo2W3p2uxNlO7JqLfq6L0lPUkVXvvGciQ+IXZxVOHsV
yta5Y/Tvzh5SfuGfcBkL7FN1rr+H0hDfJ0S2hBJG0nErljlsfnlNuRKmTP4t+e2J6LV+meK4lDE6
rS8ITShDAj6W71kpjfsON5AFJIaf9GFSR/wq+symLyCpZ8sf8fBm5izITH70RY6Y2APIliShJi0+
ATwlm0dhiudYcy82Ett7Gul5nG60eoRdqabfOiOi6A6WorA23yO7Fn9LDaXv+rNpgdXXHsODwOB+
Zuv/S9blJ+qSftEpZhKMh1EvGLZzGF5Ta2J1/zej1Imm/q3kf5a6oOle20MFu+STLUm+nRx2mhvK
L0Ks7mXNyBAcimiuwWXqrY4LC75Z1BObA7NSMW9qqzyD1hTzDvf+6ZkEcgJ2lCEGlarXvKUSxGG2
VHPnaB15qFlrZhCfOirO3hxZT9ADH/L4kvNqSAP4GDExlsjY18FLTrgxnJkw7KIwp/W64wloNdT/
G6UIzgmMwFD/QR/k1yPLsTVLJiau5FjRORSr9KojbE8H+pCyEcznJWHuG+h9QyVFSRuBcLF6Eh/O
RSu0KlGMNw50nQxz9++OJMOctCXO6zKsP+ua6KMxsMOCDMpyxkt9E9i3VctkSc1w3QBGFQANAj+d
GVlHKsM+DASIdnjO3q1612DSDS3DMclbA9lRZ0tVh4bigPHtuQG868KIvDuWxkSVxngBDHr6N7TA
kdoebUdyMJUN9v2R5iD3+VcPR0m7K3UiWMhk17EIYRDzPAdS1K8wqz7kVNURQjbL9HXq/odMbnCV
JZpzhS85DweK7/cvJ9VtSCd7oAlT1gI1oY34G8KjqdJ8IimQM7cU8CvdMztM/5c+boBXnuF87qCr
t1kHGZWpIWdWcdGNAGupJ9LezrpYJfxgk3BXhRvBMPAfeH0crDLIn2Iuqj2XiRDOj9rwBtc82l5f
CoQ1aCmG32eXrB87/Hl9rhg2JBvea1cBl7lxLypGJ/R44hExiFeqAn0OYSWHnIdabKHDwicXyqFg
Gz/QkF8iR0gE0oOphQ+/Lti5KW5VskZjTo/UQV7h1gMOtw6hx1woiXygKbV1Y+PAuUCoN6n2juye
98EwIDyWodqyq/0DAlHjkHmx9CJPT/hxrhqK8msW/FwjmiEbr60C6GwjUzMuyzEt6NQiocI5eqei
5A1Q+zUwQUAk3dHCT0SOwKSpPtNrB4oVfJ0KmQtQ3X5tdoLH1d4GjFhyRdWB91vXiB85uIjchF6a
KQ70CxznWJQsDEap+V4nDdRGMUhL1t/XsRtG36IU57v33Nzic8vxqziPGzusDG0p8LTHmgupbFqF
mgOmBzTp5Wf5iw51Qq3cfN+7M1RNRBRBKJw16F6qb1B9KnvYA7b2k0+DXeyhh7rSEphftHPPJ1PL
20cd6wE0q/+B5dn1i/H+yp9xESOl0Md/Tsz1lP0c/ZeTBFVAeQwZbK4G0Xys74KUEh9nletNBojA
lSdasxIAgRVlVa8g8BLYqzHEI6i1MGGTDncDhrFciUF65JpyrB9kChdQTrwxHxxvirFQBsDfVtv5
mXlfHOJDCnfka3gfCRlkCYX9Q0xoCkW4zYJdNrVYVhArke9YeSTz27mz98CjHoLXNrA07HAIM7T2
NaCfHv7e4FICFfejrzyoW+tL843FMPAXPoLwYgS45dKIWoC9M1luWgywOoYP7GJM+rheYFXA3MBN
58AKfNNX5T6/CGsi9QcZ2EjcYGPwBzxigxb/bz8/cWvOLoS44FGLj2tpCwFyn7ZG1FJwr/SgQOWq
hQfZmt1/rZRwok6hyxYxn5ygNMbqTw9IU4J6Q7OHl1Z8ChV3M34PoCSSBo4c1R1LymLYnWf4ffJr
Junb81vBrIl7+SLc/pOfLHRAUQuYBvCeKuocXu4GntOX5oqEKFTy+b38mTWoJpHRPMnW6Wi8VsxT
WVb24NUPUGBqAmRjdpbBz+bsBKB0+OZiOJNPj+1oYOhJdc21b1EVNc4zEQz9xqFTLiV36C+51oEj
o/7HWj51hdwhUHCSFFeJUm52gap3PlXKBp5SNocX6eM6mRaHyX1kj4Rfcs7tlDr4jfuPMZFgOxJX
V//no4rOAYYMXkDGzqYyqQY9BMhziB30olicS4PrqY32Dnz6pCvXnAcukzcY2TYXxGPIYURZtu2M
pkVnIcUDq4i9nJY0guU79Fnek9qk88hjfh7DgEvPsqg/Wf/S85VLMnWW6+hCKirxTGqwJLto8AqW
CvdBpp6VAuBB6n7UIEfUxtFWzbAjwd6cBxtQtwrD8JtnTKQ/pzeDqDNCk6FZtOBUoyfX1OWmf23a
QYcnY4tQbyUbk+eT42HP1VKnVlc9UNGNnHuOdZE+XpU+JA5oyYx2HEY4rSFp8IApn4GHndvt0Xr0
h6WJVjQMsRzKj3PFYlOdS+6+j5HJHc7A/qsKuNtP8WIR/WO2URdqXY5h8t4RnxzFosbo6tHHCvYk
QdeCkB5hx3OjAxseU8Qp6BgfX+au8lBKiJ675TZyW7jmAlQkbeNVYz7qAT54PW6CvZO42LmBhsPQ
l2riZP7ObmGeH79WC8OH+CmLdzDpEv47EfG+gVS+0bDZ1u0yXCvettLljTsmjMVwJ5RtsYeraqWm
6IyUi1ytuAGwNo8urKk1CF9a2SnKa3/LpUijfuPq0kXqvhvfNbpXREXcsShGo6qQrsO6uknD7+a5
8Uyb+XuZe55pA3WUpdrlr13YhRjELc16kSDBABXqrfQXFqA5QJwaN6ihqe0hL+BavjyhJOj97d4/
9V39DV5R7j+ngt4gAAAH8Ai129iGOGpsUKTXy8ZAgESWeE603GAVhRsCnaLocy7NNm5coOaVC4/z
TALRMy17OLr919gxR5OwA5ALMm+85TPJxyq0HZ/U9B/dgSsMDytG5y8FQvuODkgBKpfloC1KPYGF
Ni68qo/c2+9+qpjto+5XUJOEgjDZb7K6EbnhorkC+k5iPkTsX0usaIuaVKg2SRKB+A5KYhXQNNY/
DFk4Cvcv37+TS1uQrRJv762HRAkdGzwj5UZpwBDE6sK/7ddogi6rRCqYbFKQScJZRERJED1m6T0B
PoalWLekf5FDhGNjW6PxJvB+r/9HqVUDTEimitcRqkFfFdTz9ZEAPpXKIjQVtma/kokzwY4dyF9T
PmQ8AwtagVJZz7WM1hFFByJff7yF/t7Mbxa8a7QTSkx+9PphER/DWc3a71CXUN5ulUvcwChgG/eB
BHbgsBpXloApipQvVGqMvjHe9cm5Jx4lDbmHPzuS6vRmdhzbQJfX41bwKwicSBC8Yw0neMVSPQPp
juoF0lWfGenVB67Zs3H/gDUQGJI9uk39cGlCQ31no3DfRKo7eGgw5ZOBRRzcfugwbn5itC6nyfiv
mr64NKAmGxWM3UwnZVyAQ+c8FOlWse6Mjb1zaNbtVn4EEj8+KvVvgSisRZKthkg2YnuV3Selbnix
v+em/jGCweMrwDJGvwIEHwBV7jSJeDaoPPrTqOWRp82VCcN/BTtMRk7nR+qyI+jXwLm8uKFUu/cF
15VO6YJhxAFD/442jIH5HsGSWBKzg1HRG52kGNPZ/eJhB2+h9vkPHzjWJUiPLQxzNKDfcJ8e8R9T
Xo4laKzjiIhLrqs53hmjQ8SZW64437/khB6vo6hrHavsQgJEsBFops0/TMqQqKWgERXaVVu7Tzy9
UmI0klx22vDL5jK95xJ4sNa9fsCNZXMY2f7Lf6ILDV9+M7aBzO+y7iMaYf9nyONl8xzwHPFK2AD8
H5jptDPl0cirH8SL2u4iY9yJ9I1zRTSxMQVLnlj7O26jsmeuwnyefdpzzaSS1por3+ajjj8OnIRR
H8J7Rj3WaxLqaROMO3LI+SMVs1m1Vy7Dm7rC3/jiobJu0lI7IFdRLN3HC8BMPxHQ+Fcsz28cXll7
XgRommGr/2ufBTpwxCUOiM+/41Eo5dfNVENQa8JzNartsPea0ue3UFrokzgQq68RctU3HVeE5xdj
xLakHm2tBCtovHyqDHA3uaj6Pc7wa+kcRv53QBzGj1JWhdQ3ZJqvxVD3N+N7OG1oYbUlfUVClglY
rgQtTjFYkygrJG3WxVpaAqynt+87aInZT4Y52ZXqVkt49i0V5lJc+XRHl+njvPcAhhb+RXZbmwXP
9Y4sTI91J3TgPWoaCkJJd0d0O3fU2gEwgvcnJFHgiR2GR9zTSkse1+3g3a62PRtrQYGilZZL9xXl
rI8dSEtSCMfIgkvnseM3TAQKBcWQPpwvG1ORi8CUbZrzVLVVQGn6CErKpmuE6gyreIblXLg3Ewqx
2WTPEgNTN67ZXNhanhayZsGy0fS9Tgv5Qvy7mFDGv8p37CVxo+nyskoNgWzWfEmBJq0aXi+uoj22
H6Noj0ToLE4Bn2WMSYaNQmaftF3JXcyTwCvoBGAXj2QzUGGLJ3kR2OWInW2sfu0j38iTCGlKhB77
tfR0eg5tVE+e2F3hXidkkFvXuOxJjSu5BiGARR4thOamkhrdJe8vjxAsFQ9ZB3DKVS7ZI9l/AW+V
SLs9ek9ALGmMylJVfIB0MWXXd0CnujMfu1mnYXHAU91TTIScb/XRkNXZ0APoyYShy8Q77doRbvvF
dUN0J2bNxqLcyqgP0l5Ifujcgt+3cj1rCgGL9RPFJDu8+iXneY1CiIZMcStsY4tdtmZyZpqYjyev
JRnXg5HOvsMcPQAtaVjKMpsy+kh2mZOF/6KIGNbnmadZU4MiFzqOUYzQDSfiJHiLOdoqjYbxOqP6
33j0m4fapHIbtWo2bxfh7aMo4XHmaDb0pZ4YY7S4jOH1fQvrHRHfPJgk08XDqpQFEATv1Ssm2f3l
0o6AX1IqX3PQrKPDHKm8ZkiVGPX804UpvF1b0NPWAuLIcqWNkj4LhM1eqG/unj8QVPsPEqmwFyhb
/517DUxp2jDwTfyDdbD5ih6+65JHE22LAC2RBpqAyfM8m37McEV7BKtryhCENKL/gaxLT4q/3faH
dWjH/E6gtS9qzy8Cr4iBzDz0uBGa5+PtnLC7ETRGNvqyLBKwbbmUtArUzgG3EPU8UJUxaKc4+hen
M5+9LRG/LG90vgAsRyXTynOe/DRGT365rfRUuW5FG0F6n1eQYpyN1agNI0SwzjjWkN54K4vECJKZ
b6xAXA9eLdWejHvEnw9hk3xRrDYaA08FsXifDf2U1ddwE2nu5Es28tsveYIX1UCFNUgnTYXzVpLH
6Ab5TZXEw9bMPfENzNh5T0Htm7SKvtGIffODTE29bNYyWKlRBSpOrFXV8iaAMRIDAg4zJKLU5V8U
F3MjD/IjK5zuRxH4cg/0fNDebtD3fJQm5Tz0Gcg/+jDLH4ub6wZ9dKW+8grqjioEvhYMecpE0sKf
3L77D9/R16zdtpQworQEwecUspCAbpS0iBT7PI6qW2VUsjFkUQIApFEdYGFIZuWYKAdqNvAZT0k2
oJFJuoHy1o4/yExwgy4X/4O0Qvvc9AHqHufEGJFK3I59WLQrvdu2q2tZY1pEo4p9NURT3J/Ujo4c
gAlmlVZuYIbzupGly6QnBkO3qumaHn483A4EeW9mm66Z1V+TaymDnKDEjKvzq6jDSztsoQus8Wz0
BjYYDO6dKIJaD44uMndHQ5+UmI3MRQ2lnjWyWGD4yQtaR/gOFBgHu5pM8ESC+GotyeD4W5xWo+Bg
Bwys4csxiVW8LbIm4dCkQOUBhJJk2zfLKZLU0P6BNKYgb4S7nXmVexUdgCcVEq8MBuQ9ANdhCweY
dbCTtdXQKAjrF2z/sObD0nM2Rg8/E26Dgc6zVIHX0rEVlMBtnvu4eX9TOOtt464cfq2rJdP9f6B1
zfA6FU22GfokCwApuXFNruSXmARqFaYh9rj6w/Qhkep9GgqBGXkKFkaeYI6Dvg0IhxYZNDDNCOTm
3w307nZ8wXX4CFsMKdz+adL9TG+V3LPZ5HJWrxcc3M8r6kDfIlfrL77Rdn/BsGoso4VBPdQkQNT9
kfjnl97Wp+PjLxJfCIXHrWo29fKySTQKxsrAxPskIzPYr0vbsVUsLCP4gUgqDhYCqGLLjojfjiEf
kASfu0JDkgO5KFgg3f7/Q++WcKieu6Ze5y2/s0J8RbBSODNuXwdd3qpHAOVqN3Mai8iouAM63KoL
FRpOUFDV7gKen+l36AzgNSBTJYkWfVslaQUFxz2kle7oWas9zTLbAmwkKRyHPA0hYL9HWuoFJNix
S5G9nOjJ1nrH4mBtnqS3I7mIYMslOkNbvvo3VRJC70YENxZCmoNSnXuZ7UvCfC/OB53fNFPQpA5D
sJrX3ZJDMtgwABqQzMyG21zrrehC4ZnIvkSKGEu0NDtQGOjxlGvVPs1QPVEq2qzkmWIobinkvkmR
7SqGOyDXQ4ZRR9GQnCvBhytyPvAEbN+n5SYU83R/kgBwrJnNkQhT1ddTcQLEsIhCqURoCioX5gzX
qVuldSRU9Xpo1wHPGMjI1UguLpeFWx9Lv455TMrXorfpcMQeSK9fL1KbUG5miCTfUGq5Gr5LwoPv
8XOz60KzK8IU1UyAn7JxPahPmd7sCakCgfxUnZliXIKvrVpHpZqjhnT5Ep8k6sP3jTeEoglN2oBi
1MRiiosUiQOk9pRhZfQEr1sXr15T1H+MWwabiCave0TR6o2/O/hT1N1gP3bC7iGqZoBfkMtHpA2s
QBpHzX5LjDZ86FsJ1CG7QlahDrrEujKfxdS4zi6iPDonUq0UAR5hUZNrtnpkSY4frgYOBMwP8o9k
PHw48JbRTLQdC2P+SaTrj7FVySyMXDM/mlzBjNNp8+el0wuxphFBSLLQy5WxyFY54jcS9SQqJ8tC
QBx4cnR8R/UtdYo5/6lsMHbUZnBH/Yzae6P6ctqZEitnfm8dmKxuY9NwwDxJdtfeL/2gnHHfqZDh
MqPIFXGgGmL6FPpnNY9P2YMTCGdGfbVGm84jraWydu+xv3MJbYx+I9Vi5ywNPfwU/CuMHpGKDbQs
s9EhzLqJG30Z/eiLw2+V9LvuXSmzb3crvrRQu9RQl01+J+sfDhLiA107RIqCjbNcVQXjHBmvzg4P
WVkF/68IDRkIaOMVhfMqV1TDQDWCqeU4GELl/H0SY79pFiTIDR7GEXznnf9wsRr6yBasj/XsR+4b
6RCiApULJoh1hbZbC97/guQT3s4f+mHa4KTcckh6iJH9pywbLdpqCsL6s9GdPpnAt0fBuy0E1aAC
Q+zt5PS+HRWIhAxTuYRA/piNmnxkcJnwRQdF9O6W7Mb+MiK326Civ6kl1Ydp01xjMt5h0hXhCPuQ
cALhl6YahRzDylIaKQ+CFg/IS8Lh6zsjWLGfLjz6eMhV3ouG5eTzIVyGzSfLQXazRGX8P+G2Hz1B
/wW5/VBCTMlDQRs5IO2+tWgnlVI9TUKEdxiUgIOwBVYsk00hjJiz4aeNms470oEbSIHqRVJsvEYR
N+1cyJfJMu/9EX6hG9JYGVUIQPu9fGwLBFI9JY1gHS7G8+W5dzoaIgQID6rjjK2vWi7/u9RgkS7M
gJ+xcI3MYzHahArjsTImO2rcir55dbnA0CpEH42d8GgeNOqn1YERgKG1ZCFZu2o+NIMcGwxQk7rB
5QFGO2Euf+Da6reVQTQGmCA7Yxbd4usor5U5vtXjPyFIBgreQ6FU5CrTl7i0lCED4zmZ13ogc3rr
cIYh7TBxuLVZcF3ioEFCsE9FPFOv2d/Xs5YJNnHmWnF0ouVZ261QIhDqzzh5CJAznQ8TH5m7ML6Z
FFYloN47GRffjojYJT+L0LC5973ebOnyrHB96Kgjom4iL2sHqpZjMApBafcH+5SpYFrzAU/Cko+6
F9HfJ1w9ChiZEA6fmvNPL2P75g8jz75QJcl2Unhh6zo9D4T5NcxA4d3dQz975sDLXW7CUJlbaoLq
WY1E7qp/vuG2qjoxOYAkFEUcpsYwX+Yh6tpBpVU8BDC2dVBN9NV8hs/KPZluM9XqwuKdg143depZ
I5O55YlpTI0ah7v58A8f04OrIHFpoFy2QWhG3lbdQ02MchDIZ74FY7j1BSNhOMlDt9WtopKHgqHE
7Uaj0/RDxMfgMuBpY2lhPWs+y+B0c7eXW8DuLV/4OUQV3P7o3PHVboiHz5NE1eZ3t203Y/KPsUl1
cPRY1+rpthtNusHgPO57fRQnZ3FqvkF3txSelW2XMirdxA5fDHLsga7FQ+WlvuUOuRf5D3VMq7xE
s7Ny8g76myuLfe5R5AL2r+zqEgBPrSUtJ3w5wqyto9s0lZdOkqMTrwINouDcwIoxoNwNPRt08pSa
X2IwNLhE0kAC5viKrVJOjs/L3or1YLGjARD3DmiSwKIpb3GMt14xelnHy/KTvz5dA+m/8sksLAM/
FIC/BgW5mbDcsvOv+UYwWy4wjrO2Uh2VRN+hRR6/ylB8VVPeGNyT5KSF3kpj6JVllsqaNIbonTwz
WpV3rnqmmFKTYs/PR0/WnkqTYLJSG4mmelIZuqFpu8nthos0mHp4opsOEr0c9Z/3Z+IaI8iEAHGJ
QSNiXWYB96TedqHwvNIB+4g+yUbuyK3Ig2QBoR4pQO2RTPqjI3kdfYKZmJ1MjlrBxoum8hwy/x4K
kswxUt8iZSwLmVJn8E4DwOQZ4XcikH7EibDc0T2CEwXZRVetM8IxG7b6XehyYC9XeeajODlRPgHL
iRfy8xceDQHxwWvz7K72C3r3fs+qF9PVbB0qHEsNPSY7V87i/x+z8POyYDI0R/RJEJ/deXidSU6C
nHvzofNFtdYqMZl4QF0wkixk1PXn8QA2olA04A2wAj8MZaga/2DHsYk7+W+gMZldoK1s1BWMru65
FBtRiNeeq1zkUjJyNhixtQV87ZoK8MCNcUSRXYGCPeBo8bMSr5OP6wkeU/KrQQWBIBPFdhVYGBGl
tcTD02mwfJZWkJgFCx+R/2Uy3OfAx/W+/KmswZjhlQGgOVezLpiKf2WU9OqN97i6NOmoEZPgxuDY
08fgxZ8RHx1+mXLd5/+uBx+6cSRxU7YTNpATnLJL9qHuFROOxwOt9jLZvfyBZYAp+Swg6yA1k8hh
24LNI6QESdMga7spqS1K3ibq9YCPvfI8ElSNB6zJoMM/MwsmNsXAL7zQamnwv2VmGpoHEuQbU0U/
JhloyRcdHJqdjRjUZe0wLPkfRaeqdta+T3XdHw0328pkCSPv+HwStjxeEzfUZ0tc8VWYla+GO0aT
MxbBgmP5TcSvzecuHK0EIMGqqFnleGRC8kIFpJrjhdDaWGpLmhlliFboh2NT540UyO9L7+Iy/+5m
If81l8fUsm8VTj3U1f9XiiuWZwrP4KF4/z8KFatK9vPCDeshrwOTyGAcU+7Vspr/BJ1vsyoqsd1K
IySWok6Dv/5ybjfWg69vWGM6ScSo8ws/ayP57kR1PIhCVbWIiQws7rfts0nueO7UqQZ7DD2YQvr0
olQO5UlyIyA0WII2yZQp6ED+HC6dcoeQ10r5uUglTJePbv3YyG+xcxrtMUVklilvXeO5GO1RbDTe
Ttm5j9+JJQGA1yrQindHJWYLfFgXdG388ANfvURVF5Nv+6jgU7bTKc/I7nF6iZft7mCWJlOm8UPl
/FWKFT0LExt5/2qPs0TnWGWNPGwWsivGU5lmoKgfRetSGpZ2Yor9vJx2DXuRDsCn97FXXiH/79J9
6w0tqPDg2XpyN4OB50VoWVSZA0Uytz8VZ0Brb+/gMBN5YiIPqxCfJxEBaOH6Hi7KSAoWgEjiDlFM
tFeQB0ZmPhjLN34QB5it4VEAoZ0ddMozk2cYSWYTacTTzXwR9yCdB3B90Dy924WnP+ES67tgUnm2
ng4ZcQs1o4jKR+7bWrP3PIJXCsSh2dHvBd7Z7lDH5nYV7vqpxSFT57THnKDHoxK3QzguzF5qjLoc
Ycgag9I6Agfety7yxaxTu1lMs9MRQf+A6RIJvPPL3R1wHgFS7ntLECER8eaJP7EqJ1599hkC6m64
tqGisnQjnaOk6H4EJD2Gk8ipzTkQp3RTh8bB2KtM9d+emLCbBwbRSyglwRaVAKZrvo4WkO/mvdiq
IBsa/fj36H9glpnyFAM4bEPPUleQr1m3e4ug4N2Katge3sKrq9wBSgcxHVFt6QPBpTKe1zEh58Jh
mMlLtmLnuykIime+XK7x43alC4c5cbNP4AiLSnYQ1OBZpQlcUPQy4XrmnPYhZ5pj5XCbKFXnRAkg
NnE4k76LcIJ+UDQxA38ClCZ2VstKuxg7E6vZfyGIMweerJuWZp9etsMUeu14yIMbosVzmmqXsJl7
jZKraOz8CG6hT44l2rs6OKdzIs1GWdBFk6hTpYteEa6E89saCFP2C4oZf2i+uAZZY30sYPjM/q32
bB/gWZJYxxXdv5jwAuIpshHx0ph1/ycheZpRBLuKtfkHKC9RwHBqamtbGC0y9kro3Yf6OUZYMspG
RYjMz9DPKbSCsi4N1q5zh1lV6Ii+A0voWg9yJyXgtUQ55B987jM/ZlhGXHCfRcxnoaZ0mfrB6JHi
iQtmp5oXIxAxM+DkLWTCS7WilPb/QuGMH7kH0HtDX3Xvd2a8uIWC7VO9Xr27ESdCw/TIffzt6aOy
C+lH4+aD7If4NeUSbbN1TCvAQmM37NVoNKIJhdCPowvhnSjTXULPMH2gmziILoPDIlmLWWs04wZY
OchKRcXmtYuIBHjji3pLylgdzSclcwoGJDmumzxuLBsBJvQ9E8hW+tPczVkTNmWAB2/Qky/7TmWM
FeBPwGcKe/1PWQtU+d6Xe3PDcSaZmbpkyBwe0iPWfIDsWBqXLjFG2jqrmJfWH4eEZ4MhCZ0X0tIH
QI1VR/r0cSs89pPJeJRBG1pthgdMaSckFcNXd2t3GkUj8jr25kBvR4DdyLreDkfnmFEJsBEfUrCW
Ak/xd1ChLdjC8MAUFyAJGkDbT9pagMiOVDv8tUXGgvPFIwcrxwbZPtyX43Fsp1a6TC060hv8MnBj
6I2wlhFX7flFGRCxfUY6uloz21uKCoBHYZzdFBLDpQ5hbI46i3zyrD2vySjFNW7MG/1MqELNRUUY
jAB2I+zQehrRq2FjyF/DJRTwnxSVA6+d/iGqM9SzltsT861scTmGMeppReQllE0KyTixcBOYIw/5
+xL2clOMdfMkzCo/8NvesrWX6nr5Jl2urwCzzUtmUVJPUCa+jSzoo9oPODgqBU36h0NMDSUYExTj
UtVK9z7e00LosNJi28EjBfO94l3gBmJQ0eG8lDJdiJrx0XWQzvG1LtTxitxmXiv9nJqsnk0HAusw
+EslO+BQCC+E0V9v+DQgNm8jL3fF1+W/JYf0PNdBZyikdPahTfkMUTw426zN8I2nAks8WYzIn8Q0
on+SZJkzqBRJa59cWSjng59TSeHGWa/tl/GRdEW4uYHTqOZVX6pBO5Tp5xJZM/9JVFN5usyVTNH0
2mHc2Z2WsDgnKfCsn7fsikJ1oEJ8FItgxolci5/dG1O2XWpxM/4LRSPTM/13Qw7Nk4CXwCwoHahW
HNOSgwlYu78+59M07Dtk9/TVUWgMNiiksVwSDJJUpR0buOqxmpB8/ScUCRXYUbYhb+JyKoy2ts0M
z5JlYSRuUXYy61p0CahYMHYIULeJrO4ONShgF2QBjMgVdIxGYji52zHaH7Ryiz4V9h6VmVbZ4wEy
sVvSWmH7owt6mBcDQ0O6obP8N3NgQmnSNCXTbmxzmXesILlI7l+W807+/FENidfj/MCKcumvE6lo
Uq2l8UjL3mDjRb4LPjNCKsNWmae845LtJWqh+P6mBQ9xkOnIJdWDT77AjnJeGy5KsZx0eoJXOlQF
QTeUkNhFCEZcdwuR+zgeJF6kDQLSOIKpkRUP6hrNhZjw+V6TGlQ1Pt96WUVX/QdrHYpe2NPlEMk2
BfTZ5KO6bOjHATNlM7ZeVRI6nppDuBwjPBflkNlflNr1N45T8ATiHw0O4BKWYxqa6/0a8fvBBtGq
gzzlCcgwSUeD5byGBXkF+d8FXSEXCAKzaeQIA4+lwrcSkvAGLR53iQHUiUICg3KwRYp8qaTlo52z
apb09m3iMg5NKwbu6zlwuTbpoFZzcfAJZSr1iOo6ZTbqG0TitOiOGRm0fe4hGqw0xMhuDzbcKwkV
tNFmNMJd9Ck01DZ5qN5LhClNHRto0iydLWokSgutuq4tO+CYbM9OfTi+BwJku+3WwTm4kEFbZZgX
z313HeY+YH9QaFoNQrbb8RZeQmvo4gODsydtkJjTZHoLvBOIg8uqM5HMlV7+VyIJUG8f7SoyJ/xp
/I51fBvW9OkWzJY0oRQAY9BVQvTKYmCnSM+Fxwz/aqhtom11PdhZs1cL5eFHlTVa1jhTn39b0fK8
5HQFzAYPxc3YwN5g0aDR8Ixa2IcjI4S+jJHz34y42ax0C0u1gdwrTeCi1jR54MTrcGQRWVP3gm1u
7lw+BpiRwKEtYaTYr4P5VhssirnNdaO1ziXjGyU/o10XOEbyfUQzAuwWN/UvKQSdAyhKIKUtJB0h
tWNl8YwiOvoDfbcX/JGKtuUG0QCkigzBaTy+5ZUSDDCde5QGcin7DGkVgZoft/6SbocHblq+XWz6
OmZxtwsNLUmIs4k+k6gZC6H5Tw97/ikWiNvG5TPalUgHdJ1UgeEwhgbTMCqwi6L+vvYAfo2axQ3f
YF4YJPYkrKVsRElni+k8zAUiN3rqIerbOEFahHXy8s/Ktzp6PF8eoPUc8XTk1BH9Lw5fsiUrp7bo
r2TjfwS5AWO8jqh5nIrOjXt8y0hSb0cdbn2SxBnoAwKLKnN8YhMKAa4R0E86ArMTve2b+qmOkAE+
oEifHQOyNJr9KWX3bBI0+Kpx66cj6o1g0nn+dQm7QM6NIt1IlANXBuH+VWAfK8jXUJfTz5hsTPil
49+cUgVAKmfcpt6vMYoIGp0651tA4ZmvBdEiJfOQLaN3W1dzQbGGdRgUKJPt72WQeIvC117cxmip
PV5Q0F3dVQ+pwtcB8XQRcnjcDc2LU+d96FzxDJAHvF/YJHHKk0O2ztk9qXndrg27fv49+DDNHmax
rwBsA55fQf/L10hw2824/o1YtSpHbad5fY402uezmxYFiDI4ko3xyTYpBzT+yg0KWYH8MIicRc9T
O7GksyNHiDz337m894rLRiDdZAmfFa/uKlSxB9B225voX7vh8bkH509o/egqci23Q+8pOlejfK5d
3B51maVOyGNkOubFf9xB+1800wvCZ0gYtQpGc1YlSr8BKJ7PB15bQLa4DpPt1G0MtPeO/YlfCl8w
SmWRDrIu+c4QOJfZrvH28SiEizH3ZPsUcsJgMgu7XUfVh2Dn3ajPfG9Jm/FlXTl3MamB52uazgZp
hKPUWHvTz9Wka2y8S7h6lHHhhebsM044M1ePnTL4sIrNzZBVNVHq8ohRQISIMd8Do/V0Be+HPF36
gAz0yTamCPtiKd/Sn/g91F8Fn/rE4spatq1Lr93uJWkesbOWBfgjg62pHnKvJb9Ktji+lax5ekzp
9zEULlqaLyxLgqSVawHmS5XbyOnljz4h/jZaiXivviFSflYQkV0X154Z49ail3gwO/mmEMh9rzUm
dMLaQAWF9xkqS3FRBp/TvDvbxaX/v2XNWP+Qa2IlsRTeLuPc3EuLemDhw8Mx3NxQn/gCqVZGtLFo
k2K5R9z6Vy8z0HftF9+GLjRGy+ou06AIOB0DsnJoizPbLuk4h4Y485jqOwAwygxMHClPeqbOTc8S
sF+HPM0dbs/jwQ82l3+ihVd3XSPwjOV3XL6bzj2dEPCcseJjP9u32f5BBICOaTtcOuGMM0eTHKMx
u2BScmdJxdPnLM3Z+TjYTjkdR++qNKKBUpchBbzMtuYZuGjJcAY0cKC4dhdELEwEFs6GxctEFTtM
aqSvtrsatOQejcRerQmlQ/P9PiYTFSANLvON/tXyI2WBgs/9JI/x2nxO0C66xJvOJZWU+Z6p9RGs
V7TuRGFtPqNd3b79Tezy7mBu0xPRqDDpffBfbvPjtq7MXKLVyTPf/Ephn3tczA0Yrdhq/xCjVnuI
5AKsPxjCSyK9Ozo7g/kdMlCbZPIr98VQ7BMwnh+x7vcEokaQF/wY2gzpdNW9BFWyuB1hcyvWEnXm
w6Gk5vAbWetFbFUjT+vh3FXHWK9bpoJsp9QK/oeR2jXcerb77Tal5ovsk2DnTltJG69rXCfS1ll1
GBlt9V48/I0+2yS+0RiqI4X/V5U4z28xX6JEH7p3iEy6eLR0/tv42+EKl5gXybMUlYGvezGHgYfX
2gjkvR6qrz0VM9lYtNZQkr+ImnFQm0B60gowD7++/jwTBaKMYGA54//yqgEH/+EuvwMWnX/fdnip
0OrE2BvYvpXRcPpgkmMUQ7/uCacza56ZkgJokyCNaXcxa8YirDbi6RYQxvoeivztY0+9RjxMDhAp
t8IMDFHZU6QruboVjXH5fF5eS2r0WiFiXuH0+jEgPHmJXJcDBDm/bQRTjaY8ZcQR7MATH5sWZ5kY
3tth15ejQbzZFG3N8fQMSwBVM/pnF8/tqA4gxxtRl33kNVh3gk/tGJwKtpfUh46pOd7T3448Y34i
ghl/tedBWxxehVLNlQXo8rGQhcLuLaoDwtz07IeNpoYo7EYJdZ+3/qyA7M6c/IN1HxXb9y4AQtpa
jVLR/qDPXYFI0uA3Ggew8qk8KoBUvE/AM6HJKOuE/daAbpCAXH6mq1ZgMk8FJPwLg9Jr7BTZT5/4
Bu3QOWhns0osErpv9jmiDl12G7XoVgG5CAVFX7RVUm8BkbtHQ026XiVwaMl4S85fzZqUwF5dnZVy
IkE64WB/9m2KeXiRJnc3EanT32HS4ygAlIwQden5qMc0rfoe18icaneQuSnB2rH5HfguIcPS+nqT
IzjZqHkk8Zh/UIxHtLssiqNIbbYoXjK0GbHmDMy+UaNG/ezGlVbNHBZ0U9K8FqLCRZEx8SKt1mOI
TvkDzJyzlxsPAxDlsFl6MH7V+L0Qk6ir1CgXJ9ud3F9UA8+nYUPlZYgAMsaeXhTkzg69MqtUFl6B
J2VsAZciVHwbmX+4pT3KbuGBDrhSV3Yn1rpe64w+K6wNmVuj6tHx8zkk4n8ZiLznMyg4kawiyHTl
CBbLDi+wv5qButRvMWJ4/AYah6tBSjBRRI432AsF+FqzbZdictymQgGcgTCDEiwlKUIMIcwyUSGX
gRNJTdQ5DUUO5WmhhOjpE9qC6Ttu/gl1YlLpKtjtheG8dH8SoMPPFRRLO7yHNyCYI/E8iYiB/9CR
5Pgv5YXbnxwsdkKc4oiNny6Yhsc0SzhxWP4mSSvZyrDoCuJHhRzMjQsD5NnBxbwQMRkqQD5hq1Va
hbsDAIqy7Vdt3hMMD3INx0XQtwmsHLOTGVAvq9LUatE30jixgdcQzSAuAdepP6yvZsduHPTcXexn
oScWOFXMzHU3m+Z4/xldorYqk7h8aDz6zTnJ5/t2Hk9Lj5n2AtP43TI4HgfsxJXMSMHV81vUXM8n
yzeG5eZcWFqGv1v3JjjfwfzJymJOgM0dJTIC8r64uE2OUPf+6btAovK3kU4bGTwa/ody9o3yUCnB
Nhml0MSjq95sYun/F5DfJQ0NVadXfpED+KZ8FaH6eJb1f0nDMbhn8DeSVTMc7JzbB+cVpeZUa91c
gdE9+cteYz393N8ZiWBSbJfz9Y6xxDgybhjGx2O5Y4/JwavaXQKO7jx2roCMpGkLnWEM7RnbF8ey
6d9OtIW6nUEinMQDuWdb89M9D1wswMbAHXKvjNBQzv/db+RtLWbz2Q6KfMw619H2D9VQZo20kRHr
mnGvHkdpcJM2hFZvKaSdwnP8XbdJV61PbyoWmpyguRjHqLqIlUeTDBO52/5O5AE0YCCj9B3q71Be
uzyweh9iGv6usrfk7Snj6TifzJchdOHxqnXm+jRfQcfgJerY2MxPcMfbtiu1Nz1cNXG2IK8XgJlD
TQMYWent0Y/Z5jbNvDfgQljMLX+OX/NG07cGjCh99z4J1N/G+gK0yPE8IJNKqabS8L7Eff4pjKG0
fa9SMyd4EiRCO8IVvj2L0BmxF95eRpqXQLpEHD/Juxk89pN9noed8XKzW+GM8cmPnEW360pCpqey
n3I+I3vcCuVNOu9kixJ3IcyA54TuEFIRJn5D0cbkf8KUsn3bS9oNByX6D6JAPmBK+b8U7ir1WjIR
kmu8WM2JircLnKdoLNFc8RJKhvHgBV2TMHyRMsK32fNPXagey/pYqUxBwM7HRQsENe92qKKKxQNC
v7cyeNF5rB6PHrPttcIL0dcOkWDQZHL1ntWNCnIlZYMTv0PrWOMqQpiMcgFNo51m3s9YuLte/k1T
fJqak/LGAjk1E5NXYTKYBS4IHxC0LSy8RciXj7Ycn+an9gnWU1B2GncFhxUgGVwIYLuJjR0sbnL3
j1x5izFlc5zjpI+TNxcXtlx6AOywxH5t9UR5SKzTQyiN2cR3eqPenEtw2wnnnY3ezQWyCjtXEGTI
Icu7n0KACnah39dFmXvk/tFtI10H+pzLSfsQcXtDmhgg/04pmzqEh0IUTZNwXnj1iEzpjeaxBo5/
rymRcUaR5A4GhY/q8GfGdjp55u/0c/BV6d3cKz7iwIF6FJa4qBcxAncdCxQY8xTeK+OQ0Wb5idgj
TMmn9jKaLu2vqJi4ETcqo968p37xmQdQ72Ohj6wHDQET5tST6WdgxhYD2VrNxBXfq470pambWR6+
O8/8aHTjkx55yQDH6FakufUvwJmtNGfXLJ4aW3cJGwndhoiIRladqdc7xO3yQACFQNvEDD4W3ZLx
eVqV2e4F3osyvGZwC2jioHeeSHaU5twhZa1O8wThnyXW8BletvvmJHh3ExQeWIigFTAPQ0p75+w2
xh+xhxwjn0XQc+3/buFDJ1Wgv3JCAettKC0YH5GVf2AgaDTA2pEgs/jNCBVCW4xOysZZ/QAmvc09
FMFG1Uxgp9tWNR247nZCQJrL1yRBpZ1Gh5qbK2xTUqtZU6SUZKItrphcmjPR+SP2bPaD8ixRnyxq
/azgs9tqrirchGaIfwAuefFbGnHWugx3Sn2UvY+0FLKzT0Cc5F+nKkhSbvA5+ZdqkcNlytheM9ey
3sbma9E+Bw+2xzu3MUOEMUKmNnMjr/I0H9cp5LT1gW0OhWNjPSPa3+NalWN7TBDXV4dVsSUZpVrt
Jp9gTnqgNWtKDv895aeVs0sUEHU4VrwyXsij1nKmhY1gBX00M+irVPdwjdlqg3s9K9JvqJDJNUOL
4vKoug22PXqGonahsXooSDI1cQ/7MZjMWF9YQxU+cYsZGmGQVkc5EV5KsI3+AUUcA/VmD7zyqyNA
XuVNkBsfHRi5sOBYw8Quk13OoJY5r7v4TL4P29sLpKh8EWyWbbofWpzEiTRqzZslfcAdBYhmu29E
z3w4LDmbLHr/YJDBACFoQU3jbfVFj71qxiIEfqp+ame+73/i5x2SYxZunzBOxhzzG1USdOCvejK8
zCLMaBc/9eC3CxtGnEXlY/i4VJu6bV1NYKHeaJWHIz5q1MQYgPSRZEYjJnc+bFqoewhCdEbmXNtC
Po1DqNU19TfCxEC0GqvGm3Qe3Rgs2Je+Qfl8m7CYmeXz32pKiuXfLJ6M7OP3C7/eTuhXN+BiHgfs
2PlRD1sqj3b33VCOmYiLf/Byb0Yj0EYHM7YS5Ue91LOwO6fI+2uSHaHaha1Dy7tSWGimfzPIbZuM
eKIUwEbs0VV6Cb2YDWhummUqexr1vcyN3riaWBLnoC7e6CmQsUrJQrIVqKlRvemWyp1lGlETbSrg
UXY6lJXVSmTKqzjLZ+cnQQSOHiHLoDZL7XvU3zWFaUVQ/PnwQEmnElCZbJKLy/cM7jdNRVk+upd3
bcXGRTSSCTs/nv/1wDh18+gZ26IDFOCDhuHDBQdnFfCkMsoB249kKRCPUYC4RgZnWSNbAknKkBAe
28Din5QR/uYNIdSYUtN4afX5c623t1GlYaX846PvqZxKjUYpJvtj9sHuXzOGCSOzsnNkRbr9+BDD
hXpmU6PRNLep0I6loWIyR6VDgN6ObsWRigEXO0ithL3R5o81I0XonUTeMIr/ruKREN8HNvSYpCcd
204HA3paiVUVRjtqQLISBr/igzcgKVp9vmnj8XHXFu+lmzwK7Or2ATnt6FIn7RebAvTOKiRDJ1Tu
xqxAsev5RRAuvg0R1lhp0Cj2KJUiTKIXdxLbcZW4kS8eewIdGw5Y7RsYZhvhK12Gfv/Isqq0boBB
1fSmY4NTMHpoXkcp1GQI5NA91mgGCXnhIPRYkMYWBxwFjf58K/X4motEUkw8K2jUxGJOL/McyMMk
xXhqUvH1z9YptKcUvy5ljCiTPoEk80hZvV0POrgjkERCNfUfdWoARwcKBKM+MdaK9U4ZuTtvdsXD
6/piG9KUj/511BJbo5A/ALOxBR5UvlDeMcHQcGjhYjKBKVaXasjhCyq60WHNl9sjwWZp4zL/XwE+
98N1aCJ+rLaG1+B85I9Zv8idjf7hG+0bSfgT2h4xo/DcRJ7AZJ2m3CjnZEoC87LKdBUDH/vDHIWB
fhUzcLTLoAWfuocRtdxExIdD/c5K3Uh9y1vy1pwtk+Vr4lV6k9LlClkUTzGPcgVAgbO4O1WfZa1/
xJvwYDxOfOhNXZtGHXqSlBG5xMHKQX1bJCfVMrUmLUC8kXj/RUZQXF0zYNIWxf7gRwHSgvIWafb6
19WWUusBPvyNqgjCVB5lF35e5COvOT5F5dE7q7XSFPKUJVhpUdh34ZM8uEKFS4fCWW/V+Y8jHgOu
4YZgBZxndkUR4xukcS0ldkf+jCgiFeXn1FBtcT4Jn4lrY6XGSI7BVwyTldcf77TW4e+jqO+u1sRH
x+KU9UKPt2ECSj0/QIVLg4HuhUyP4wGo+A9/P3dPU2xVQo5R3IrYMdXWtOFKbc9/aSTwcPXITuzn
5bhZygMvVFPnWnQwg+LlROxkYn6xdec+JqfU5tSpn2N7SUABKD3hVQVw260UleidyY7lNB964deD
uzUpedD+E/Qj83vMTRXJSZhQbwZMDyNauvaz2bWFFQImQSfsc2rcZYH3GDDq16eY6SgGajipsPFw
GkpAYQdYtKQg5rUmCN37/Cq8SpzH9SuHdW5ADGiVm9GAtnl2P4mWA2v8TdM4QmXLF71r2p0npFZX
8dNavGzTp0WNDJf60oxotbGE94z0SbV8FaN48YOBbULEXikoMxJWWBAtgyjoJEy39OFWQqP+CD5d
Fw6ZXQgMFdMMEVdnZF3edHWUiIFu8LAYo3p4AgzDub3n6FVRhdJ85vj+SE2HGC6srRtcYgWKIadk
pH1MKTyubiYUrwJSKzYDja6bnAFvKJ7WUgD9TiLfABtY1gpwRL6pDXW4epHJUe2+jzl1GlvCqGeN
Te715pUSbZi/kzOuCPr73pf5L6JGkzHYf6nWrSY3vtvlCEs41uqmhz9IBgQeSQshz3SjHvTUJRhq
Msf2zs6q1WOZU3ikCYht7qhUdrrUh1gs0DhJz0XUkSMA4BmYTiZ0qCyHWeM0q1JMLbnCgUzck4Zg
s5b0PS+tywsqeylNHgypkfMAc4aN8cIbFCZ5pK2lXHy/E0MB/V9Q6ie0HWEnbE/sJPXpseFiqsDi
kyDvtNt2yQPd+LOxnvXvrCJ3A2HIb92bQHHhhrQtD9pHNzi7nQAvbryoH4pUixtJWUCjcREwwdAD
R+qjW1dFBit6yuyIylOqD4RrepFFPq8sHqNHQrgrjrulylwywvWobK2UPUXaZTt4CjQ9KO9DYBdD
umTKOEiop09Gl/0HJJVxSbNySEVqJafZ7g8UZyWwqhJQqgmLrRdIj0k0YCO/vqcPo0GNXDJUFlEJ
je0wnKdSGJcVC7s0V9QYoO0LBwDEuvlr8lvhX6qfj26jOz7B5Kk79pmCPJqf/ylEznhfdG2tit8a
I5nOJhQyVYcNYUpEZ0cU8nzRxWX9+ZAKvOmeOLo9Vmw2dJhdR9VEpUfN3kmm9B3DJwPb0j2LQ0Pf
fucb9FMma6lWHlr/IhQOhvfu0nFQJtDZE/zUoeMFVpimlPnW122B40iXK5CMWX8TIZXm+kjzCxhK
b1c0/KZrl8hwtdgEqt9YUz1ETg8vvY3xSB6M8/VBUgow5SjCPMOgzLQcZaubSgoVfCEW4fibG4bB
8JFk0NaSQvC2oO/qmZJ4jXAGR92+p37ykB3Tqik2tw9nVFnPKfu9q2Ig802qfWEclecuajPB1+Yb
nm8HGeYmC9VNXgKDptiuRDnXlm0BSAoDbGo49jBP95vnqHF9ogGATy52i1ptteGTv5ZW2guy3e1g
J9vhyC5Ldhj0SCOYwyD+6SCTAWHbYcdzipeI8DUxJQOXs3vx2rWl/+PaucBW0mDM+PJA84Ea2JUC
cx6GXqz4BkjI9ggYBpqGiw956tpuuH8hw/eFGWDq6bvofOCf0QnK6I2GREtgLkXnnfq/aXvgiUCt
I71wMRiAfsYqOsqqb3rm6FE5LqC0K7vpZfWCFTTOGLOf2VAwn8eRr7MvC0VTOA1yFg4Tztzd7X0B
N0w92x3On1s8GwwGZUbIubOsXvcdSuwuPVYNZ6ErSsyteurreXsZ9VVrmiJY0eHRUCpbW/6IJhmD
SpsnBXswLRfRDpYtkONUenShviIRckUWlt9TTYO5xWHSbF7IIXDNO97jWU4rMC0zhkDgiSuQeJH5
2THDOysWObPrSBDQ+27uSHpGs0pt4AzQLObZKEEbWXcXuAQdAj9GLYZUVCmrLd1KwivC2sjqMoHU
+GYrrqo0IK0y0oBzybQudrvxkCwt3VlhDdNvLNiFaBoBfYx+8PNpqdpyna0Fu+FtJfCQ6Cmgf+T8
2ygSWnZAl7me5jNfK3Qrryaah6x325LqUuKdr/0hPXXI2DBHA2/rJZZLQl4aoOEKKaW4+iuWZVaD
6sLDg/aQf2gtX2PSES3s+1APsIst6aSvFmjZBjJzmwG5tN/W2utLchWbH6bPPCGNe+scO6kiBk/x
XNVirMmtdZ+kKjOHcWTMuLOL3DSKTCprAOtlDWibJLA39c0AIx0lZJNixDzFOf+DgGtwNWM4LDNG
lgjSAa4z3bgW23a+MprbZ6eGR5FI3qvSYwWYINDTQ+k47Q1acKfgXHyRRB4/qqbLiINiBaPHKjfc
jzL2CiyrIa/cUeSc+D8LDtcttbwyAGBSNNJFoL9l9DK6GMeQtQasa6Hhk765HZu6AReuZBj25ftG
I+IANIutneukIEIOoE3eo8bjQcbGN215EP5n7MwrIygIAMIL0Ns/+f42nJ+QGdvRXLGc6UBHSksl
TZQdOSdqIUNomPZdqQaRXThQxs1uS8oCrQ16pRIg+ZZkD9giXHRHH0axMYcoCVM+QjlPwblwx3W+
YPJCG67WYaTC092QAqUSqPeukSLZRCh6t4DgQqIc3cEIXypFt7yp95g/FqYPdf4It4OEfcvNIxcf
h8hVAxYOSWqiSMj4sotLBgiJswO41yyTouSPhGwlZXkmPY+Fq2kOIpwDsV1jvQZIoILFnPsWQ6C+
SsDy0G8/bm4V86v3dvc/QybSKu4i9vtV+k8O2mVESxt+lKLGXrMbzB7AtIajQeNAGS8GvZXE9INj
n4l/Pu35ax4UMHKI4og3PGqFtfRmJl/gbRVZmZ2CuvcyqK5cIVFMHeP0j4uAM2Fqk2FxSNUV0LSs
piAEMQ85XxRA01SN5C3yXy5IIXSvnSjvmkDicy7jqb8Qe6qaD4KGxzoEne5YK17b4+FLsqn63bM9
L/joji9QhdwICiYI/7ew02p7/fmfFU9Sd2YIOctL2VKagvfY8mi4EvsEXy9CfmADxVXHpFW0h+1g
aRQhcstGHE1I4zWyB9wOzOHHHu1weIUpiLUxvgPFWf+Fxe3csH2u6oWOhDxrrJUbcdn4DdZ1bh9h
Ex2KNPzSmhI2GPSkqbFDGe9mtIwCMExncBDkEGNshwDtWjxNRym63DsG/BZ+TEBu8KgvJOmO2gSk
YDxH6G074Vvrkf0aVDtiVCrOS7+R1CDFCKWmgsNq3NbI2610Z5BNlA61FWnynlkzqfEB9PWSyYm2
YEb2bEWC+yDn3S4di/UAXC4vBSethBex5v0uMyYp8ZjMxCpHIeBbszTuARr168h/N+cGIiOgGlzE
191ny0pVIynjp7dhTQJreNE25R5FN6NwqcBZFnKM7xnVg96YyTKgpaRRxQawZYts0ZBmA6bAUxWK
ivMzUGtGlXbkLXBKZDf4GzlVoUk26cWued1vCiFQY1bD0GUbr+9iZkiuNJUToov91FjuC6QXyLhn
nP+Ny1T63u0FmBoQPMbBxEPM0/twCYfRHxIou9+KXxs2mDrgsE4+/dgKLQuNtpuGq0gFs1D1WDox
IBzx481/bHDvpo8mjTDwUqJCv27UTDqXxQFHJwmmRVxXExdQCkaxtxlxi2B1GRX+LxkQ1Oe8NDHs
km82hLCrcuGs6deHug0s3hSZas8KyQiQT2yiYS2IZq0gzj+34CvOzUCgF99PZxq6oSLqMUjCP8AZ
BIZxfr5V1Uf98Y3eFK93oThnbBEAs5cUhkPkCcbWWzMWExL1dBRYoWW5C8o61/oqjwRUzWrSfhnK
fxc/5lEOAnKqONvGRV7DpzfRpQTMaWNcYIwMJLfeh2BkRWIhcBGOL/29Gq+VtZNDfSpxIx/yAkgu
A9xQV6V5i39ysOwu0DD1i99tytELlKJp0r0ouXsr7xo9zoo6jbtDNzxCc6ZNyEJ1FO3ebK9H9t36
lFi9N57bha89KS1MaAo5Flu8wz9+wdcm4SVewa0c629yz5J0o6mE64F4aZE+dk0YiMmVVGaHmnJm
Jxx/OvvdUsNRuWqV6sos+gKeDX00J9ul5un784xwfa9J2da3AGgWIlJa130dKXzVim+3QLT1fqOn
6XaXGv/YybAxW6nfSntmyCcpU0psPCxvwYL6Si0lohh11uWhtie6e/ge665cPhU/lIyvfz3Z66+z
fdryH5JxFwXlKSvQDo7PGlWksidJFgD15MdWePQpXLSWw+/Bhj2xS7BzYtU5FU+CxnTT4MN00c0H
PB46srdbGMfMvhXEduwaHmZJn4pz0jhHaDiAVY0tSFPAWvCXLdArzG+DYvYEbkP8jMUf6veuuZ4n
A5lQrrSeGDGjJ8h9nZl0o/YChIbuIQoSPdaJRxmHEwlxBNeU+lETIrsP2dxmOlvWor1h6rNkRbWM
3ArZYB6yRZ+4MBwF1VJTv28AlW+sQDrkqqfEtL5aCTFY7hZUDgZ9KuMFiHg8EIPpoQO4i6ynGHOt
Ei9AqLZ43OkUrMW4qKrcx4nkEZaX0tqWCW7MLCAOCo7WUF6+alKWUtmhEpK4TfYUYfl+nHPKo9O5
ANk6/xSC1V7L9sB4LqeYAPlN/zNkHfXHqZpx1oId2no8ratDV0w+RicH9f2cG/jHDq0wEMLZPJam
BRn7uF67oAq1GwGfFbjKUma3eUR95SPHrM6urOzuHiHv4qEcroyzQT/Gimwb8YxyIKVjn7M7SCzZ
tD3NR1ymcCbOARA6+Zyr71+GnjLw0nlZ0y69IYv504HZQAJwFhrFYATXmmTEcTAmthesA2oEZG3i
DwpRk5+TvPkAJlC0Sk0O2OibzXZIi6MeFiRAVk6DlCXcO6FyL16N7Kq6M/kUKYsWzigjHSgrksZc
h/+WHK6FeJsomQAX7e+JicAVvoFM8W6j+Zbza2cJwX0WwSsuAv7oJdDMraynwbUonUo4haDjpROJ
mL9G4sVw4hG3HBk2GnJpBpeXySi6sZNCztA5u+5rT+65ZIU1waoQrbmupUFQfJOm5C5Xl0/FPGmN
pD12NvyMndDvpxjLF1DYH6kETdJvszrodAJHJI3TB4HhSW4b7kW46wpYzwATSI045o2PWFifDtEe
96xPUgd3rmnUlaqdQni3TQs4/aWEPl6MLSEwiZ7P35tNYZKn78ux9Ko+87g/HNMBE/OdzN9ZyRq2
xlYQ4LNeLRteT26JmSDGQYRajMFjzW9SCDDF0wB5mGJbeOR0ilY0Mxwg4oMADs3K+q4mUxprRkMI
X1EiOF5zDmLbahVYmDsWJnUpUT04mSnuQXlf7k8bBuZDC284Lz3CfLMyHz4+xk9mg/I3ReipuKKg
B3F1XhCPJDrfS413mU5l06Ust5EmXXwFQ6fEzMHG5TxtHamgznZRqBQKSD5nfud4ln0l6HieaGPA
17v/Qe4tefMcGo5/TMJLM3wypb/zDqwvMo5X+sZ6nj8t938legjgC+PL8GF5Tt/G8PW4+xGtrYfn
pFQcIEwj4qQ2CrxrLQs7MOW/6BFgWZcjHosxrqoD4Z5QAeRj0ivgyC3dCri95YTS3xUz7Q0Xc7UL
QD8UQw8pUwpcRLM7sGHQuTIfjid1RfZldhCboo5a6Q/E/810mcccxubRWMZjXmRxtDwbrUs0Ol82
zIxurM8iL/xm+IbWa1tvQQzSVGO7IBrollAWckC/zAfJM431p+aly1cEcraxZvspgi181scPviW/
hP/jJkk5lLmHjKxEB9Cpee3cOOw51u9n+X/WqhVNaF+DLYJeAFG4WQYzAnh1U0QZApSoUGxbgpA4
vb2I7gx3UBgHxLcq7udxKxZra0Y1OGj6DZ+lWESB9xii7VmKXFavXC4t4oI06m8D/b27HeMCvJ40
b7UODT+WI2/4k3OztIY5OWvUWkK42npCNFxKpiCEdwZ1ywt8LdGtnmbRQ3Edh0YDtBDE8xajYelK
EuKIf+lu2BPWqCJ09Fp4H7NuH8Q1kzLx7f9QSE8vuCgtUTim53ms/2y5ln5pLJYw9rQ1gTxckdP/
N64w9bx8eGETtzzZuOn/M4R55+lH2Mt3jGVw6wq85FFXvJrkV9Ohz82OZZFtgrPWlMRoy1D/lg27
3WdVNOoKidpbeysV+EV1BGb90hnFjN34adNA4igjVLnP07guvI8eUHiJFEvLfEAh8rblA12vh/xW
RXqjAo0wOYLmP/wHZMf4bzqgsYduaFDgEYcprca28buF25+dCNGsOFPCSwdSBAN9vWT4wQ2dVEBD
2ExtzymmOpwAxtJUNVDwQWPzKANAgvOSdSqq3498hBWP74TbIq81Xj8uh/0DYduMicJqyFF221Fk
gSn6oMramVFcT93ViIH4e5RoBxGjxSVtlVbd139ZOBQvUwUo6K6aqddWqzdyFmJHJt3mUDKHbS2e
WcVXDiS2cweBVlxZCE26JY8Vq/w/MlRChKvhB34AgzEVp3vbPiFwYL2mgyAvTzs+6XDgH4+Ka+ba
+IVpamnjPCAl4N7w0jBRPobQv5rvQ3LQD2OOwwOvPIq6pXRQPRQ2JvHYggm7MOWzJBJbBfimotNN
4DWkFRQM6CVZmaw3P7EDzushv/SmidmOxvI0jCpnGEWl2B5TVnCntz/U/2S6bD4c0XtoQk2kvGxr
elTydWjC6kryNgAcvDsQMa+ZgIqBGuoMZZgT8HSCzzsH1k+qGj7T0Cu7kqN8pGB3CSzysp+bKMC/
tNU90RytweiwWjSjjAbUSF8VBaBbFsq3xQvEJPqhpcpwumC5CyVOfgdjz7SPKixwxX2R2vCy8FIF
gdzodiz1nGWm0HEPEKxS0pW7TsbQFhuc1zgKH2kap5k4q4IV0QfkdRlDKMhOrrd7TQdXW57Zt3Go
fgz7Mv50uKj8tnOFPPdESSxBrLKxfb/kVLVkp7ruy4URtLTp7KOlbOPXJiInTyRMD5IvbnNaHlWp
ROQipCD1AGcCvNQxgI8Hv+YkKnJXRGSFYppyHU5YgM1puccjOl4Y6MsD7cc1XdLOcILWyQaSXIKE
r90Pts6XHyGJgsAYVDRoSHkhbyvayLx3uSEQ1mpbgttqXLoBgug5aAUBaFnBy8qxo+OszHnC+A7T
LUh4MWUiltNKhNR9a04bSVHLFpJEXdJ6wVSxFfP60w8RVoD2liLE670amB7RCItbutsq/npDaXRY
Q1cTX7RWKc2skc3pDFXR5nDF/AFm2VscyKPclCdMdcHzx+FtZruvYJkYxYYRQ8vSQoDM+8nkC64T
FQu9/C8vQbRkY9BFK85S64ZOTpqYYLBDWxctVnaTBNZMOwFcQITD1JbhNe2fy6sPsw7f6mU0bh0G
+08BFyfROitNdJ1cIBEzOB9yGXS1cInvnFy0IsCh87RAB/tiPHBWYqoHTOJmLaXbmtQOeoq7HZW8
ZKnJKE5gy/m+mSnupUPfu86lLgPbc7LWsqLTZNHJsyO9jv2SkxGcmL0B6oPi/onicNBMgN9PMY1N
iHhkTuGSNREIKYdYaGa15lwA7Suyd0XOl5Nzbeew1lgOCZzAiUmbBP6NCHHp06hS9GZMsycOlHcO
4IJu5tbqn1b6mBGLGu//YlVggw8Kx1dRYgLhB3Q2O3Fw3SAoA9GEvqWeT0qAYOBYoetlDZ+g2opJ
XdYXFrjqfXOj2J+knTGMiz5CJKvTeVZLEpjO8FAOQV/VrAgEQFDDFOOd/2gvHy8xUxytyBv+eMWO
yH37fmtpLVcd/ww68fcLLmn3EZ+3b2lUmmkwM6JwZuadRmntriNQSnaeu9jrqAf9KnU10MdNaqpd
h1Ya4U1uRETXYWF2GvKvSEfS85Wyzd9QZy7ojDyJqQgjAQHWtr9bAX6tdKd8CK0fY2Izyt/BXRL7
5jLwuyFN5Qwu6v7WirKI2O/4RZ0EHLrT2+Mzswg0v+gTKBrUkVMJf1kvHbSYz3Ied3rHrnMUb1HU
u8AGwcNpfR1ohRLd/xa/9retCmsIvpumpDR0bq1PtfCooNTglUB5NQoYx1iyOKxZvR1CDX7mURB5
lCTioj6POgNECWhs6EYgFG7t4DKEfQediM1QZz1A1oFDK8dFmXbckdeR49TaO31/Hi8M9hijOwPW
Bhj0M7P9J7Aou6qIrjfVQxphM6P1JBjPkNaqgYhKJ4B+jp8XsWbOKV5Sc6/D3Hr8SQ7ljoQg7vna
Uk3Z4SI0nDWdEtkNNW0/ECEZcViRT+qmbVrJI1QJsq/jX7iXIuscL3Zelk2r4yLxbkz4M1ZTlqvJ
lTFn5D+5vTKcPRU38fa12vy2UPydZVpUAcIamjMk/eRUyqy3Pm6obm7PQ1B51qipeV1T/B5Hzr0C
IvopQ5kOEOqd0iKKizMo8Ol2vKKfdUcAxl95oVkEyHZpw/qtq1dHm0H+kQZqIN4bwFhBK469iuGD
+tH4U1EYxnYnA8LN53U3g12uN2mpgf7bTFbcJxvZKy5pkCpp130ByrN340lrui9pf7yY1aED2mPb
xgPUaTl7VMhzK/JTSCnkK8HZclNMClxNE/Labuv6W2j16+HqcVWZEIRQZDgW3Fq30tHPkNBYNHQQ
JwjzoNPvgglJUHrcHMw74cV76x9YV5Ymgey+rw2UmeCKug7I9SwyuoDO/EwhOO3G0ZZ4KZpbmHvu
fP7zR+KZBJrasPyFQ2HGKhSJHwYLDeOnmWHFN6rmXph/dmF1aesWt49zc7LlktP2UP7QogqQvTCh
G6uUDrA5YBIu7nRmtOGUoqxTmpGDuZ1HDJz+ikIL5Zs/HFoJgY2tsKZzN3/CI5jRxAfA9UvjiBNh
A9WJI0NjSnBhTZ+tRS3xA/cOZ0tutx8RHYlikIYBaVWKB184XwY9FID3J2ds7gZ5iACcZITWtc5w
KKzY0O1hxzaDkBZoJ2x+YsrEaNFX+0Y6GITh/ptiVC5r65M7NI9VxfsLPYzBIjZLHoLBVuPQ3o3M
f/ViByTwKAx6bHmAm2n4ySWFZgl7jEAPGCOG2gO0aDLxtSFC/NQCm7uZGS8lS7FiZPLsKI+3lLgb
iNLn7Uc/fsmczKCnzAn3H7P37Bt6y+uimeh4gqGoJXvU5nkUJi8EiiKigGdPPtPMFW0cn+Ky2tUf
+Li4Rapna3Ae9GoEQwsv3Kjsv3yPoKBEeSWnqzpB2hK62toIrYOKtURUeSH206wdpPT7B1D2Lhko
VAUBG+qBZgI9Qs9di6t5TUAjFLXAVHazpY1/6dN5H6JXpWB0XznLG+J72PnOn+vJIacE4+FPr+9S
Lc8G0Q9I9UB7VaXjq9Dad6DHZzH0USb8lxuboTR/TsLf7Ji9OczeHh9HtyRM1PrpAhXKVccj9r96
nPJpBtahTgV59XYGIC6BOExroZyvwjrp5VQ3nPZQeKC1CuxU0SIgKgoEjmBNpCNbVms4fu7y5esM
ot3IE4l4ukBMZlUnrNa1maaOLX2I9VkL/aRHkJ241G13Z41CDzA6AvjLctk77qIVmH29TjJMYqru
ebs7nwGOtTBiW/pbrukKNZIKTcpiCbpCmOhE2fT1EkJYSvUm1LXKxVwKuUI9dln8OjlbVmBJgogW
AuyJE0pCZjLCrYiLy0FeI0Q/yuUyIClQV7FtbF/Rkcuzas3CoBsXfACq4/RnfDctoU1wuCW8Q/OV
ZolphqG2MqM2B1E+Q2dsE8GR4aGl2J1FkP2+ijhPMHMilOXIFNbLh3oP8whOPMsoiV+BGQs09hUW
0AIKl8WT0OSOpAJJsg/fXxJjK+/pc+drqV1Yn0fSceNojwiYG9DqnKR+nhAAbNY1E+FPko+eJ/iX
0qukwEuZUsfw8p+0f/J7lcq93xJn4GlNY7DZDTMn/Cc957bRbQvoNhjnojIuFC9/PpVzVJeZSocw
bjx7sRZtd2svPFCidUIe5Hm5Zjf5FM9l6eQME/AZec3v5vmVWxQNTKyjbcz4W5jvAEoAqqK0lxys
mJrXGH9CoZzwUBjW3uBABFxy2h4pFPLAG5k3qk6Hc9v7QmOVHWTjRL/EpM8PlUwRjClGViNJaayd
uzEeWaRFQbdIeTtelrXa/Qx2WJtzLKs10xGuKempEnRAs6etfJp1w71oF6WQdAWamZV/055TKixn
PxZSRBwMnMS/vqzj/3s34tKHQYUzkUGlYLG2yUjor6mVpSEm+GJ+o2+14DxY5I0RKLim0My/eddB
1BKg7o0MBgw5Jgtd34frROVYmQV61hwO4wUygPwpz1srAVqNbIeMfYZpP1FaMssTqpK11F9ilcOZ
Q93ymMrFcUp92kuyD7U4ZVdoEFMLPw8VIUVwJJBlJYFBRittSIYGA4DYQZGAQyLJVLS6uB+9nGf0
dvUyrgnC3d1oLsMT590sCuLIDoqzbD3Ui047u16TvXoDbNgiBapYT+QD8O3hVNLWMfPxGDXwcTkh
uL9GJRvmB+T2oMg0AlWhU9cG1rbNyA/uZE/6l2uhuHg3lg/4jE27TTVI2wYh0RIxjtdac1dxfNIZ
8odvTuXqdl0NWmSwXo9y7SdG7jnxEn2qHvjXZwaAE+JIfSnU3/eruwhuWHyXsfiUnCHrXkv0t7nG
xrkBflZHvA67d6CWbWIrVoXYCDSca3RcAMGhNZzYPK8cIJUfVpRms5v35Oe/G2qELJGaky6xhcQ8
/hhbOplHD04foNPRsfhVw2oU97pizQrOCr+VcEz9mriLrEfE7SGwskh0hvAZPtSWHSVF0JvQ5qVt
AX8/AyspAZjo9tjJ+YRhwp9IUYNDJneDIrIducHthu0ftoGVh28Rt7kEJ81Y6eUTUp4HThMndI1T
3Uozy+AGJGF1MybOLrq0UJACCM1Otwcpe1qnfQnFdXWbjP3rg6zNMIb61FB5bKIUIhiyt5qFusv6
/l1F0RVqvSNCxVb87o5o04RrzqHQfZlalkhts7DfsXJUFI08Xn1HNKqdkgSMqxD05HqyanqvGF/m
PhSkD0LrBmI8Ayg0R0MaGCkio0ZEjzuBXscfgH4BOBba5ru/dgB53hwnf55zXRS6007CtLR8JsbO
nhUt5FV4Nh+9t0LnaaH+MXA/GnA5Z79EIHxTaM87JVcY2B7t2x5SJKsfVd5VGz+se0GqZx5hyNTB
zUx24d4/gkDURD9RVGL6g79P9B9WoqwG1S/HtsMnqg8K2/ICLxLmW2Q15W0W0Tcp0p9SGKIfb4/+
XlacPB2HCAZheMzmdpfUwCnAPg5vu6S2FqxAGEo1Tvws0WvDJk6XGLLZKOrnZMdhGVDoG4B5237H
cpFV9TuizZRhZes9JEXXZpbr/oBZnRemKXWaoMRHUY8qYmFpDTOKev8YwOqZDWwyqZBW0WfR0q40
ShbEsoNz49yXoCp7jUGU60k+BnE9hcefgMXciqWV9UQ68CWiDDSncFQGOJPRPbk7FQ88MLsP+pCJ
ONvAnV1MX8P8pR0smy6xgUnrn82pTZcRXu+E8nDLzQw5mpyXglfLO0L2x3TcQSfBQdNzDDb3O+x9
xmE2M+soAshVEmPuYq63Jm2DROf/37WKOvc065gaRg2Er9pcI4Vp2b6QnFfRvPphb2QwMbDmjR72
Ad8E3lYpUF5ENO44TLVuXzELkWk225F5zSujcm7+Q4APzT/YiCW/J6UsZliQkCaVaunw/Hiq4pzP
NlqYPUUZ+ETTIBPAR/TbkjtN4IQ9kVb3RnnYTxqoF+YqR2xzqKMyzUCrVmCxenK1644uC/scPyck
t6MtrGZq6e/YdhnDhksYbKqCYzQerOjvp6SLa0MaBWdjEBlu+xxxCaqXp/EKRh767Wo9R9heXp/z
0zuFSTQle7gFLWLN7D6ZD9yih3QN1P+MektqEO4eLg8EKy6wMV+uQJ2UTzDdV8O6Suq7pPPGsE1s
6yOS6vZm5w9GFY71EdZaT44WB5A6IBsMwg62Qm+5w/8Y+UXVU4fkLL1UdRNNbW+0LN53K2vyUQ2m
KpXABxmG00uNByOYSewFqgl2v6jHD7OxGKIGnIP79C+j1av5x/Nt0uIDlFuyolnWIOEFT85t9EP0
2hvTBBrTmeJA3eEf9WfwpDDiqbnGLaO6BA7mW/sp81SeH8EYJetas2zTVrcX+rBL5V9/W5rDTz5w
RmYoVyyvTs+2olH8xHkzyYkH7bk8V/jB6ClkAagq1yhwgki/qK4+2wAxvZ0M3iGV3ncr+4zwMmit
1IAhdHzw6nQ1mI53B1lNtcrjnjzVGJAx+57jqCUILtWe5757s3RR+zOkvlsRSyRZ1NV5IGLzpY84
iSm/yXUL5WPZFbcralfWtNzrm4BHMhC/91R8tcNLxM/TIjvuL7F/zfK5lnngfOgNeKd7uaAEN8nV
jS5KaXSWyvnuMR64KrTM8tQGJibl6GbdwdNIqBmrG/Sv6+iNdIos+v7MHitISlm15a9vIklxhVvi
kAPqvK8apuxb/XNXyYqBeoIMs+x6A03kazMrtIWVLacePXB7rbBvBLN++OC3Ax5kkyF/hCQS4IYW
dy/xWQ3rlD1+8wTK5VeSDXI0TyKhH2Rn15ga2vQ1qbTYLxoC7szriahn57u+B5I4Jk5UCqXkP5rt
SulwbS5EyqHjflzm41NY3bsfhJfLfYnXlhCkWexC6uVKITlaa0VFBN8I0KF1rHbv9DArA3vz89tE
V/AuAH9mZOC8NmyQuqrptHUIfVvCbs58Ic3BmBspZlqs4X1d533VDVpN6dTOXPXlZi4Rw7jumUIh
1snOxy5VSJpA0vapD2OZ2aDrc0V9ZhbmKb0iEoI4+5hHYMluIgq8EcZW4cWmzJMcQl9xoUTlokYr
/mgEjVnbBKNHm88MXYvup+QKc6rbO90/1Yep5r51VoLfYTLVi8T5CCCcFkk6zUoLzrQ3sn7J0ySQ
UREYKOeSUEGYoK0oE1z1IB1UIwiJAxvJPPgN0xXuG2hzQsDv2tGQyH+uwvrVgd8y46WfHRO3OCMZ
JGf0gLcIzAM1nzy2Zquntdr1sfST9okSJUlgJcQDHFZOzJqLCTpMQi5CA6QOMM6Qd6+kFS0/A8JP
W7cmlQOo0KXHqOAj8xe9DwxCZxsBHaa7EX51AN1TGDM7u4f+teCS15yTmLVXhAsLupE0lD27z0F7
qBO4UPhNAPX2ytcWO/oJrkyWxfqGppAw71Hkajcm50k7f6suZzY6hxBXuAejU7kkHqkVzFYH9eiI
9OjGU6I/LhSBk0qNmNSu8qZ6SuplH4qGjRse0IHPWV4nffz+El0iaXjF77h2aiJPeL28BHxtSVC5
MU+oPezbhvpJnVAATf3slRumvCUYFmVQfMt2J+lSJTfWUWArmXMShBp3HotYZJP0Cpne5urdTJ/g
COOpsW0Jdc4GcDtd1uxZuW5VI6ICa/WSplnWoMzdgLWODC1QwHBOZQBoOPmFYpQyyUyayaK2GOnW
7Rkvh9S8d1PsXy0wDk5lJq9/L1JLZaQVNjmwH8KWfNmur2Bec3+1RI5ciJjYFXw9qoGh4jnog1tP
OO0nzClOeF1LWpDHN6XWY/yIyygJDanihe0uTSgE38tl6vfEbW5AhILoBtUD3RWsJBNGpNYOyJJG
G5P5vWYnLb5n+OW6++cS6HoItjlKLhefz413pLkH5BfOG4U0ClQV+dt5rA1xCh+sA1CRCs7PmXRQ
1dipqA7X5vOz8dXFlgLCm1mA4ES04YAGYnUAjwb50v77ERrlPeDJ9h7kXRhJBdtbkWBFN7vCCmL/
wKSd4zaUXPdGaZHUlSqkUHYycz10j3xaF1cBAwxBgJjmRgv4eIFjNGruwIm+s1ksJzAsoT4md5C2
SEBBRJ8ld19fM1OjV3SVsVmbdQYuW8SllW6+2ihW7dFaLMIO9mIdI7dhusCiGYv+K0c5mGR1mwW4
tkgJxbOn+J4afK11NbBudqSsrQ4ObgSCtEn7hnPPaCqaMmGQLmop3zQKxdbSC5mU8YdsqZ7q9Gxj
2s1YMxa2D5eoXV6tk39lnazPRU6R71xNIFp7NYmqXnrlo4oK8M85RbgvfIcuf2vDpao63kQsfazp
U475yMMkTCwOmAaJIJtiK2IEzoH1gvrix2MEDXzCM057X3eeIUuD4O+ocQPsZjj+wjG0wELfreGu
xiknKp406BzoZS6GFS0EVL0+bgf+Rr9OTAykFtphHF+q1QWhrUGKJamDYKWjskOhqRAVlTeDMzh+
/Y9c/aWc9ZDiEyQr+moGX8Iy7hxlo3srvegGrX51m2czogtKndscZw+mVsFIyvqNOmRHseH/wP/i
rdfXPJxHh8mmvRLHhKeG/RAe8OIEYI8TiyyuoGjhvt3s68fhFDjPpcwCGzVMpUnTD2gglak9SDCo
vtvC52JFJAoLYoyjuFcaG7vg6c2yWN0rVSQDKQ/42ayD6pyfo0gQ8d3c2WchEkNN3nxJ4I9jok4Z
zKFJdmlBZGtdyR9oNaYsrRJcjxdGTWE5zSKSP8l48ExWRAD11OPmgILVPekCqWwxaye2Dh5D2PaA
4wmbPRC2hAeTsStL5xMnnEb7pwk+2f8r8rxWo4owNDsN/8Wv/mQBv2G1nWgRAlBh3dVagjNCpalE
IVSKTpy+VdpAJr9teVGmsyKD0xkb5b9pmfU/1PUOEZ6wGKOpQ4WsjSYncJc06C6NdDxHowB7KCZ3
QiRjoYRCCcS0QHA7r4mFXKCwXysgp2t8Szz1ULClYcZn2OnpZqr4DouilfATxiZSkIDZ0vFR5N5U
S2ECyHxM2szAvE5VUpGfxaiOk65m71mmJLUBV7Dxegc82zMiCH48/oqKL4v7vIcDfloR1EWiF4/P
VYuPKeBoBQLBDDiHZzRrdRkLXkjITev12NLfi4SNpdCZvVtnMr4HUEEO6IGRC+6ojldPqzM8lzX2
GZ8WHF8lMm5YvVhRmLisXaAawD8Dg+bm/Dt/4xfFkA5fS8xz+agc1Nj/YuOz67RDQaCh28PjYaon
xuocl0VpZv7eTHUHTo7ay87fABiShlX5FYVMiU0OB9w/hhvg4gG72kMZ0DqPOnpZ0Slco7viOzTY
dXccBd8n2voa+3ITv6nEf7Y5MN1oTeML4wfPoDJzjIBoMByDUTfIp0Endnot2CKoYpbwSirfdGUG
r/JXq39SBrXIAxJiuhXAnRGEhgq5E4Eox+9E7x9/L/ckxtwwE6+KNm0tLXDL5N8MPDVMNSOqJXFE
s/qQs2apxiH742+1WPCpZJ1dZxDAJCrgkLMAPALWxTPIqv+6Y8/njrQRQ4R/L87Ro8G0m84SSMmJ
1b1hZO1P3aoCqtpk33h2yDiu3tXiDikun8ThJiV8nZX76/2KndSkXhOwSKtI5C4+Z+7O823mcrRv
KGOsgLVaoiUI17LwMQe0Ltvd9V3OvLjXcZA3rvY+AjjUIYWHZSOb0LXKDUemdiDt/LwGnD97YVH6
VdkFGwbt2uwb7BObIvwnBa/l/uCL27DOzlP7YeBg5qa4KR8kjqleDbltuqKjdKbWOrX4Zm7sq+NU
Xl/MNarQ0rWBxc6GB5zYJF2sHS0ZnedZK9nruE5Z/2mjm5dyKkrW8eFSfozpX7n8eM3Pv/O7Q45g
dwhe7VORSKYbkTkEqB7WrYObFQNUWAfxXoNC6TQLBt6918ow7aqhzi2ClMedpt0im5KVIUvF10mK
k5VHpfx+y2lbOSoaHkAeO/b0e0oU5uhx2h1ZrSvHXsB07rccEdvfslzRis/b20bBwLFjlx9Cg5yK
6UUyqHcmYnyBNH4Ynr8COUQk5oaUbdwHi7q2+M2JoZsWwFuIHWbUMMylYfMN/8CJqgLVbbWTqlYW
x8oSkaNTOca7JTkV6Lj7eJ9FT42terE7iUmyG4H5mhqAaP+tN3NIoxNK6Qtm9JN09dzbigcHrmxP
ZxudNZQ2GCmMaFlE3Bf3GywcUd2WH4isWVLMcNm1cM+tb3L4fzjVoRnfj/5mtc6CXiwn0u0F5UN2
LJVGSFzQtfM4wzJCGrDwyNw1xBKXFS5Xxh/L/rp5y3MXaivA4UfDZVFxiuT8RqSQ+3R78z3J1yUt
ZI8l45YpIVFtJsu20V0F1hqC4TSXl4SFD+A+RUeN/3Jc5pLqTR38rrFY1spSqcNeyrNAKrzPctpO
fFpFT/RmS0utz5QMJIpfIKXk7qsFOB2Z7l9Zo+bU7Q5KBad6OyRbZvjLnsN5HbVAF1YyFpi7rIq2
2F9lOgR07abRK5T4AVwrT3Wi/RDr7i4qr6VvyGlD+9ItXKff0zMr3jK55wB2LzAsksClqdw0mI1m
pIdBAB6brMN7CvqLxCLUijaiU/WWF6naz1AbfF78TSoXYerQC2Iikqee/u9bmVdiWSMZJvUe1/pL
iRlwAPwEjk7ohMKMQE0nJW5uzptkRNCivDihMbYB0yqToQIQlRQsIBX+ztmGOhs7jpJyoMyiYa5D
QxT9F9IbWh0HVhDiRAwvTWfKIcaEDZF2twMuQlBCch6qwQm+c4Ihml2S1BdeWqi/axV77gz1kYZZ
+auIFwI0UQQxxOieWYvo1D3cqmZGyQbXL9t90OTFIj51YU/wB8cL0y7tAswUv9fjcS7+B38DXjyh
TP+sTew/GM2SRUIT9joyDCgexjsgy7uEWbeCj6CGmOW3XP90x2Rd131i/XqH7ivDdwcvyAykk8n+
Ns7DTesevgEtLijr+26zDtyNSAPOh+v5usyBYDEidHVYe+pteEGW7DaGXcidRw9BS5RT2+KbWbxb
5A8V5+E0xivJfvToe4hN93wt8PVJkktO5a+XuEZ7ssb4dsJi7hhRS3vmnqump1dLsyCZqIL4oG4e
snx6AKHBvheJdehGMaFrmDZfFQg9rXrNx1npBAROairz20tgIudowyOV4j+8JSbiS5D2ueQkqECY
ZUlkreYARz9hua6CKOUQiKioAovV2I+lhU8ueQdwv4Bk1JbhQW8szBPn6EoCDqEGE6EZW1uvzNg3
EwtxjxGEUJnvIaZDb5ixmhhJCppQh8KgLkAV5dplVDiBUdSXTY+MHmuJkFW5pcYAeIQqjPUkgqtF
JR8Vx8ngTuvevzLdLzS9hjN8mU9WFHjyV0l37kcoM4kjRzm+McmHGqKvhjS4OzQAcayZhWRDoI4f
jy8IFEmKlA1zAddkGpQBW/fbDsM+QIOWvDFt0/rIT5SqJFYsdCIEBNg4NzElqW1mYavyhyOrJQTI
X9/Y2c6Z6ivVfu9NbyM/y7no0hv2m105SA1tdg55vVRgKK5YFCGLGE4SwKHSMRAXe59oveCv3CVV
oIbAWHkJCqm8NEn+xWgXoz4UTkYOtmbas5mZmIJShfcUIkSP7cta1+PMIlblDA22Z+qfJryglilI
tfUVU8WFPxl7SmFKWJlmWNf1PiYu9XBevGzxdIIoW/J0qInt7WyIhPyvlUiYPWNkXc2QNGGHq+jz
PFuysEA5EkNuwsIVD17k2xogQauYFADeoDufvHrzKzV7MdLcxoVfrIdvmTH2VE4xdpfL1aUBXn62
k2oXLa2poTt1J6y76llfg6pJRJrBVv0jmvfmUlLzJnY9+jWJgH+2DF8vOJOkLYsZ/VEhlravTt+g
+VnYIszlLWLzc+xfgRTr0+/ULjiTfbOg6ROQNRpbBmouKO/0dJgBuUpwtFUJawVvUWpajQf4Zl4B
wemFplaP8w/h9Ikw6iIY0rIGHKO+yU3EqWrIVNpv9SSP3D5vqOFZIFOfilz6HBVYaEVKVP153nBD
cZo/cenKMUw5AgHNchdThj5+HfF53FFv1xcD5U/eSpr7DXkE7AoGwWW2rPSLVQ+WHfVBMNeFvvWy
Jws/YM5eMHTDftqQyt/h7neAri4FGvlO5VyJb/Ne9i1OU4fXdcndCxwzNGEAyycrERgfJ0jkLkBV
9cu5d9H4BWuoOOxZgIpORmdGNB1u8FUHh3R8L2v/NNUZbOxCWRKeAI98f7XYqvmmtQ8gih3kyzbh
v7yCeiSIX53K+R/SGcAG5jFPcTjnzHPAWa4Q8PfGa8qHO0Fe3LuZiEyx6AsJc1b53YxUNT5veNW+
eJyiBLdbQ6vKvSG3bgZuL8/Wzw2UkVk81w/pQA4IPqf4FGqbvrzENhRt1UtjX1sfEtMm1J9I9i5v
RMXwZSrzJPtTU4vTvBPYFmJXAwGkao1PfLTDmM45ReY+zs3TL+9FdKIsBTobkJaFYAbo3CKxIetz
WfPz6Kd3GXiXYmrfJCYEJ6V52ax0K4eSeteNKdHDEgD4K1t98za8VjkSMvHHFJe0VS6/8O0d7rAP
zsBYdq8yA77LnLK2Ptiz2rWvzR1qXLLJdBDfGO9N5HJrhJQjoObVuoZYlSjtG7pXb+l4bhvTJN0a
kzkxlM0Jz7GVGyukJMdn8rvE6gAOZTP4HHAvYV7kU1jh82ZP3Qp9yfdtpTfU/csfmRYfT7KdkxjP
RXJ+MUf8WmgYSRKhicITa0IzWeCpDyn1iBMkaVyoEh95S2pZ7C34wsl6r6MQSTWqiC2Y1vRYWhYx
QJQ5paEh3KN1qDzgQEVtoYfFSpTD3BATT0K+GfVISP8U+oqoFvVMhVdiQQgWvtQQhNAIzAA0eUN5
pGihiONhal/0FeRUwAlEebseFHKcs3nz4qB8ZtF/5Ie3QfoOmTAUvaqFJ2St6Yf1GEw925/671hG
jeXY/iCsrT2J+qrXDHtudXQP6BNDjWkEVjm1zjE5whDJqDtKLKm8qpj2QORoDQ4gEJc8eos37YLb
xQeLeoh1soVQtPb2eTkg6tAa+4xZfNzFbazliWOSJTsVKHePiBuijhZJnIi5N22kkkUl21/z2UNG
qdvHDvec6ZsiKT0/2OVz1oFhyAYMDTHB1+BfggxTtibnEsPnrjw8HrMm+w2zNTed//qQzkDLyxj2
JstJRSqx/Y2LOCkrQ8VWvKx5QNkbXmaG5SIQJZKLe0bIrtGGJ9sWjXrueUnBZ9WjGTXoCgM+vOaw
CpUy1jDpj/hQxM2iZZIX9ykQX4iygqhEJXEfXDF+mBwugmVZ326PmRs8CivZVGOR1YAu6g7X32P6
IrRduZe5gtFfA0OBqaSwgQaqR5d3algY7sPaKaYnMMviQ0hOvAQHEmzBb7m0LN3zQm2lGfZn8AYR
/vZ6shsIFQlKF3BkOLZbZ5dbI7Jt3cmsmqcvCwvG3+ybW1Xab7DQg4t3Lmoo18kOTHcd+2am749m
YPk4Frj1IOz5Yv4TCYbVAY4GVNipPnF5e0CD7H0kBo8u936iZEOa6K2tVNFrugDSBs8z4CrPPZbC
see59wn6w9twjFKF0zR7+EU6N1M5PcA7WC6EYlSWSBo5ma/CUBpGB7twSsdLYvTCDofIOCz1C7Wf
aw3tp0W1beKG1nVlppP1qrWpMr6zo/iERsMT77IZFXvrAnBNWGaUxidm+TIdSHCe6wK1o3SViSfU
6ywxE1c+zTHsauGkpsUmxZDd1n/JFkKi/uDUNc32UdXaJKL7LcJtphJuQoz/t5MlY32Jsv6VKBo4
2jEAKnVp3fcmKqqU1Zv4Gk/xntkHUIP9EUWGoJ8a4SyuNTsSuLQGBon570w0iMmS0wSmeUp+kOui
V2qz7goO5I/znTqN9aHf+4cXqvfInLtpBtzapXsynnKRWCSFmUgQCIFN9abgfP+HvWgGvr7IZU/3
X/IuE/vGpltZ/EfRqdANWh7JjNcUhkAWjXOXGsn2bKAnbOZ5jprHU7n8CWcTyyy3daTtPGwMrGgp
8wnJPebfc3I4oNdoujargQOsA8tg/0Btjzld0auUDsQDx41cTMnturKQTaoJsHkYcG/HGpq6Ccnz
qgMBkxZMeywMnrZVJN5TcmwgFI9goYYAUJ41hCZNvPk92iP8BcnohrJ5E5zFEyqcyVa6rD1Awh8F
JLRVQNbj3Hg3Wd3+tErh08qXfAAfRI9KTzr7ClGwZLNSpXS1OnV8asxgnRlgDIJypJ5jWlXFtb12
fBY3VnIk2y2hk0t7c9cClXHLEFm2h2dnuL9kPhVNazACctCACuTJMIQKy44D0kJvMUQs8RMDcZbT
Q1BDV+uCgGqayxi8rKPlnB+XD4j7fMYZNu3kNzsPsCbJGF7SDaA+BchB/hiPRyAnpl7tU3gzg15d
o7EmgSbhRm8yA4MKZuqT9OIbCQKYnlep06M/cwa2W/Zn3AJMRvqI2DhHOIJ0DFdkz6+hv8ACdSWe
oiEVuZc0Nf6SAkx6w/b1KmE+X3W3aY0FXVK8mI+TFz5qf3uIl3Ol1b65CDi+Y00kjowUVKO0I06U
KIAy/1kH2FS8Bc5O941xiSulW9KlnqZV6SL4Bh/fjHzu19XWPBrwCRwyo7gm40f2ZNU56IA+BDJH
aiBujSu1KhzT1zcgZ8g+e8QK31TmyeRuSZJVB4MFz6riXHp98AgrM35wuUoqiMpTXCjeR4gqfnj+
HauYKQkEoKaxGs9U/hM37t7Gx8Bt4j8czRiiMeUm8DW36lTU0grnj+5xYI6kgkUJtRc95ISKeqnx
oraSyHFiKNfMQxPYLnncOTk+OJPxyKeKkSxInxw0LRce9sOZKlbDF/nzMxuMf+kNj8EeldQyuXNy
4AkZbRJk+zphi3fX3nz1gpLO1gBQCd5wtzRJxh9W7lrInXlPY0ymP7hLWbWxNvUHKiyLbGoLkPrB
TAssj80VbzuGfV3RkdGSQ9WQ/XaDTSQJyidbDSyGaYh91A6bzzzzRqJxwSa5+EuBkLaVDesJIpRN
slkDzSitINQJddx4sQueZ5U53QBGGMft1+gdQYwv374VxPFVxrdbt8RGJ7ExOpNNYUDzXX0nbwA5
YiaFWv49QCjobOBx13CZZyU+Jw9MdNlNVdqjt1/7gYVSdtP/DGiALGqXHZiECDT3xNnzgS01nA8F
gmF6840UdJ6n5wDRg4F5T1EgQsQzrHu/gK8p+34Wkh0J1ehQPb84GB+A6o8u6VhkMhamg8lEdXeB
mOBjWQY/5qOG6BoplygJj8QAEOhwUEB0Wdtqozpl06dfd0466g/n/R/8yWcTDa47BG4SJXW/eZzr
KYxT+3y1q9eqf/NztU87n3fHqmK8S07ILxLPj6NFuVlF7IL6sCsgKbSmHWdiq77OA9cn0qygJV0A
pmQ4CRl9EH9ZS3/YtXRPLLWEDvgiwdLtoogc+R3E/4+Cpm/gI/o99Vr3Ii0qe1ewh+y8rrFbVYs6
qC7agDNkHRbNVGbcL3VmNLX/5DEGQK3/zouTf0rnegKNgdTfpAg6VtZ42QjxmmHjK+L69m4YdGW2
dHH/viNQ82bDR6S+vq1MnRgpNC4k0SAjk//QdRMOW7TlYe7kmX9/7eEv+eIHdYP6CbKdEMjaGdE3
Uk9upkKCzmZ5Tt6m4lPZZxkdOy7qLF8m+mcbFbR5Z/5WBmUY/SQhJq8YRUd6UGHokVT3ASEc8eVD
O+85MTrbtORUAVWjqrT77XswdZBV3kVRkt5KXBg4s6F8vflHy7y3UvlkQ9dDBCNkb7Te2WdYoZhV
zdsj73O8UaodLutp/uWV4vVJugplqxDS6RM7AxKxMsPc+ZOMawtcoH9RQkzeBvo3UBP/j+t34mDF
JkglHDOyK5/FcAAulnv1bzW1P8zJWDBlyJTmCAV8Getbj1rIv5pUdaPjehxAb9lsoeH3OyJrgmr3
Lte9EQTy3RUoxU6mPou2PlFfs736z+CEkZcqqEg4ZtWRvtnTbcpQrYTAHBvXDD6Fl0jaGKerZ5su
nBIl1Ue91ONLg8UE5+Jdvedp2IkFp+iW7LJ/sT2rySNCDhlbRxqilxVFY7H6PW4NlruLdbswArrp
wr5OEBms+83LB2jmIIFlWjT94gzXy8vEhcTKYaHcvlx11Kzn3Z69xJC/J4bha5sCRW20o7WCv8Wd
GkcasYxtqTKeOu8q2a0bsAfDSf0id9n9glbKLT+YVt5nh/nG/jBgaXe7CwZKc9jMh9xFbAgT1ezx
ICpvIuRnt/Z8QyIr5RlSA9oMx6SLyNteZHvFnIjelOlBx3gFV1mnfeSOo5ZhHzfmojJAyP7suaD8
5pcU1jzKd8hqsfXgn7C0Wz5vHinyBboNrBLdBWVft7Bn25/eLKeyderiajq7DNjbKAzk0pHtuNBS
M6MncuExk0yOmHLhOJttP3fn4TMkhCTaFBX5CP4picnQldHHub8kkJSKeKDLr4S5Cp/POIUiwxEU
MgK9ldcWqAlgAUmemPZjmiRJY/eEvRwktlpBcAd5nRx9IVIz8G1FYKmX1V+cm7h+9yjwLVXp/nLB
ddKGhzM8Bobn9Ea7vLfFXHHEGiliK87K8scfSFbBhE58DD+ffaA0BpOzlYNf1HVOkIxgOy/3526i
tsRFnXKeztNNiXeTh8m50kch/ZxewcEicaPJMf8mdG6BItabCg/f1fVASveGkOod8Itdq1Ji+BSK
11Et7o7ulbQ3MyC+PPM6bP4YmNigdW4VgiGoGuVP3xMbYYMiKqfDZDQWmd3pwr7j+IVHV+Rf/vdn
i4fLNBBZlBZJgtDh86u2V74Z0X2r/jogqsrLC4EgcSWlA9aybY0KTPIRxRLxEboh8TVJKZSXqGdy
78WZVR3T6jRxk5Ra8W81ZBKGDYyKCPe34ZlXJOFbsVr/vP0GKWFnoIrvGjm4OUy4Ty614KsaWWrU
kkihg0EMUacl9KOnyCpGGIrIwSXENxBZ0FoBP1W9+y5LxPy52A1QtUEsAKF2K62fzfvlNE9o5S23
43MvprnYlvW48D0p/bXVlB7/lBh+4N905yjerRAwxkf0F5ByJ00wk7olwvj264ECj2XF72z07oL5
g/poD4PO5P1vDU/IVhDUiwo6oVd5wqEFDTgOhIPGcJwu12BcY+fjVAFze12tFk4pWBF4dfxQA2Es
WN8CM9cLI97SylffQPUCazYuVXxILZpbuU6MR73sG1yRWm/5yP83Frz0y1B9RsWYSpmaqtT3AP0H
WdotTNgC8b4lqGL/iCSJQ96mJRnZJRDOTirwIDdXxNksQWCtpYjy4SE2nC0Wpz44UJe7TNsW4G3G
kRXqnxi0shI4VyjCuDgw0HGUlKHnJPkVUQU24Z91rJZBsNEYnd+d3T3/QJorsT5sjOmtt0938QUS
86xckhOzxKLX4t9/vELgau4aAfRIj/7xHjYKbZMGN5IfXqLyOJINz6xZBkG7AYKnTprTe+TufBgd
VgRGJv77kt2BTVRbOb6JhMgCAJ8FnOWI41+laEVJiO9+Okei1OmR5tEIaVmE/J19DuKtEE4ul7zQ
SUZLTxgvQxh1vYPBI9Wccv09cYB4si95PMB1JKhNiNhuYLJh7F8pwFluwLgoBPztjZibREkbXu1a
5s9zSw1DSiyhxgpwduk4tn9Uu3WS+ydHEYEwW2oBY3UFNxJkMVboMVaJwGZ9000wqjUKTwfogCFG
nWjcSKSeDmydrrU9jXaSjRyL9L5AMlmyw67OuHCarevcJVBU21RqC3eEMV7kpBi2hxZo40UDvNk8
zkauoaIbQWJ2KuO6z5kiLAISN+KPtwckK1UrQ3VO2YTMC2ugGE2EcL0Inc2dK/2MilrcV1VZi7Lu
joW5leoN8ayxUKoF1087YeY3YoNBl/GZZx+pMpgfyiy7uh766hj4BekfS8N3UoLBvO3xACCJdk/M
sPyv5btbrW1ko8Lm7a0g6/zcMGp/8Vq3yCLM3sYyNvg5VNshza+onjrgsmEuDVjxlAUK/z4nmXoQ
ggH1UazNSzRqbwOchTjtQra0veUbl1tghewnjBsEWtQEmE2LaVDx7c7ZspuvvZM5SIqmyBpNnEPm
9umKLRlEUcxtoO5OR223JLtfA7+GomAyvheR16OJF2PhKx0mHO0QlyCQEgaM4RKFObkSf8ffKTjR
aQpNRiD/JRJgOjLOksWeiM/4gaOw8dMtCZF24/TsFwhixugYpcKp0HAFNcXrRt4SnyiponG/G6rU
ytR1K2g8zb8kgqsr9/aWPJHMsUwRue692mxY+SzCMkvZYkzpy8lNCh68VwSvW06eLwmhw6yElv72
Cv4Qc0uxAN5V2gHOyDz3DgETZswTlxaBBUnLNIm0N2AsNL1ribGicx4pRpIHaVsJ4k6IVInozqW2
h1SAhLlZa8Zx7h1eQ9Ql7/w7KkGXzNb/S0IabZe9Je7UELBK6A8WOJrcWIoCdkC1OEbisAa0yreg
mAx+Jjlb3P8+vLQ4jOUB3BQEwZps32S1PvO3BBH/hCtq941yAuhSD4XZvhcnRiysQEF66weB5UhD
OkK6vKp+mAyZnbcjP4e4E/YHWJWyL9KpIY9axLQ02GP34XY+8mj6m1r1E5YXi7z1RlNgNXIZRN2r
zxXuC0Wh/bmnusQqb1RMDqlMsA/yGJreQKh5nyMqa+8TqBCs8HSLAWgrzt2aFwx/ANP7fVBpemZ6
Mzpb5Z3jUWhN97jmqFRLc8t/jdAhR2XL4VJ8Kdk0MUpZmjYTFaoQsuft809qTcAGyddRpU75XkkP
DDAG6LSf4BT4SOLX84oLryoMXi7FzihN94d7p69Brh9WZpGnFT0dlleuAJBYEisfoTEQIG0O3zt3
gmVjfTXSEOhJNEM9xpAcqYwCWyd2Zy7N5tiwDu3pPhtQNWtFi8OKg+J4QxjNnNXxSCFp+6BgSQsU
3x2rcSLMZMoF7/coSpA9wSV3B2mTaUKGPh5sU5mfvX0+mlaUTHXH+MW/lEuNiFIhmurROJwgGutv
koFQDkK42scZYpWThrI36ZpN0S1jXDPk4YUJr/8e7/op/UBwvl40jFt2uUXEPOfS0Wb+p4XPUEfX
gnTeDSltmOFIx8KIqeVU9A+2AAE5X+eKojvACS+9M1nriJD/ejhnFoNArOe0E/gDB13Hs+FxOYuI
QTNAAJDjXp47aSiKkdIhJPAyaL8BTRyiYr1B2xDd1sPYcP36K6/JtDuWF27wJxW0KyMzK8a+YtvR
5JgyylA8dCT5l9lDKR6uCpu+7arpG2iNuYtQ2zrlN9fRkD/2grRY4djcskD4UgEbuGJUEE+jHqFs
OCdV8VOrXyLMBgolEoTSxyEkvZFArETnxRItNqLc5aDxkzA2uYVpuEmPN9RowOkCZZIzkJXp3WtS
fB8x+EiPxugPnx5G7ntLOhyMea/F43Pp3YKMCO67QR4NccjydZPL72zMCiDwROg5G4P0FWJk9bKN
qquah7ptxrPpluVLkgo1oUhvc5Iwhe0nSH4tQ44X7TFGsWg3lktC3kSa/+8oQVxiYrVwzG6w99RD
uTiE/uIHWQKSLY9PoTR1vpuapkO8jONnoVN6lbWCVWW6gUkJl7+3Ve7J9TAs9qkxiKpB7uIOoTcT
LX65nLVZ21iQXjm78PKoWpTbOS7v2c2VjDbfN7a+E/CMn8se0EBzTKaEgG5tBMgMkeSNAzYD5bhP
PHGiZ4tColI3DOI0kBz13Saq9HwZbPEj5rVEfB+AzGfX9yQgsLYE4Op1NOTjwxPUnVkwog+TXzOo
BoqWURHSemMMGr1a91ImOtvDR2xV56pwvrzbzVP473iFnefGgfgPz+/nZU/S4HwotyXvVKs5XXwz
7mXluuFnRNSg09egomW5t4CL3D13ZeaFClAsjdPnEvzoRNk4r4ugsct1YVgEnUsZRsw3eqbnq0UO
2Q8+VzSnn40cajVYFWx1jmkbikysEL2JKsop/jGU+sivc+QLv/9gUMUXgkCOou/qsgIHoRD6aCq2
SSb7PYF7DWcgM1P186ag2OzAnqd9bBFwN/jef9agy+lXLJpeRSNwlMvrBNTUxnQYntBYyLSuhvxh
NXd60nJ2xLyhc+yxJMMedUZ0g8XfkLyRot1552DzWH4HlwsNQfq+kDOKQ9Jtg/cHJdgzz//n4JVH
7PgP0GJdYEoie9PVKxaxbSXFokMkndSry205Mxl0/xy9kUwfekVa88Ztz2VyJXStgB8rZuAbDN3x
RxP65ud9eGd34anDf0twsFHGMcBhgdcN2wAL1yJ+C6bO1iWo7YpPzaO47p58neAG3fX/MQ4+eZgC
NB2omuSMhjnd1XQddgqOTUI/sU622auP15XhXCszmMHURyFUzQyPIM4yYrfVXUlgZhZzXj8T0O7d
l/ccyy15+EZrsIfWOVWOwcxNRndkFCfAZ9x9PXNoNJqXgZKpnOw1wi/GBrpZOrtwLRc/JeagDtw3
Wy0gs/RiWBD7LMOqXDTqmv2tJDlERg/QO2756aBfU+QpcychdUalVis7t+atNe7RaktPV3YhZ5yQ
TTK8cwdxydKfx23TZL/WUmo+jQWxghdjuqJbpzBVFCi9RYkoOrbZCLf6I33JsxZVhfQRvmp+ohKi
x2P5occgk4+smJ6kEe/nCGoLJAhgetjYKbIJEAbQS/jbtC1OQvpZb1OxTONAsfh17fNrNhFDmzKA
o0s7h1zRz2ezaOoLPgzYVyf8XMENoHuPDAG2LWWgqLr5eilIOXnnkzAPOGjsqPqDxCQij+Nw6vIA
Tq6tOjcTrMinqlbbYZCujSvzy9wVdi4DFdC7q/9TQf0/Fx14wYLgGDCaah+0HTP+cy2Rqp7QFIuH
Ahs9SRJs8DfT3mi/5e7gURuTbKFdrZu5MlrwhgdkJdCZDZpShS7ONmcl8vJyICRP7tFJ9S35xpGM
h3fvxMfC05r2Ewq0N1e6QyIdiie2CD+mGvsJbruRsW7hTj5sfJMF0hlZUFBi25mYL2jrsr6yeXK+
u1F1K9vM9kfC0LreWxuc8ROvEhcl3io5QBUzRjcjpYjYLAOYgC6UGkxcaB36GpXGhV7mdt8ZIz5M
RIqFC6IR9U2wHJXYzzkCl55y1nZ6s0MhD348+GFqiV5J7oofhlnE9hGGRH6U2JKHnG+IFe9X0j3n
6FZyxSg6xp4vn2U/3l9TKjizBiwmbsp8ccIBMiNxyp6Gt0YKnZbtWbwryaw8LhvYnRMfCv9MSK1J
Zzz8lY+m7x2JvxWC3LhUIUzHjqDX6i3n27OoTYvdizQH4jqELDCeUz7AG3cT9LX85lGcMo/xcp8C
/E+toIiLz0FNXynOcPqBeYd+LeW1qFo9C7JUyZxM+rYrIpKVAa/vKmXM0nHZoW3oHicod9HJSeMf
QrO7ySh2SqIuSG6dNJGbNcpH4RLBtgmGVgietJ775eupgE5T6m/RQVosvWH1zIRm/uM8sMeEPH4v
tRuKjOUIvcd1QNWII36CHYohuzTcprktrlI2RTnF12NEN1wGWtWP76NLwOa+BW45mwiwIic9xLwN
mWL0I/KGk7Ku6YBIVmFI+SjbGa9Icmbob4xSAkNJX8yQn0Zu5SbUHbf1Mq276Nqcuvq6UoCIfogR
WiRAmKCSwIQnQjlHvBT2NG47bmnsLaNv+jDkDTdH14+C6AVA7JbISFaFch+KVwHSag0aOIAFkUrB
mVpFCwSfu6P8Fk6aFBc4UkycAZGP8FnNn+rL/YPOjMgC8/d7rJCt6B63sn7Bi7/bQXnk1hBoZlSO
LsSttfrFfpihLOJEl0oVlZKr4JVVmwuspT09xXF8rQbWO157LUKYoc+9UtRp/Ojq+7BkX5g2520t
nprWedhRS171xjasXcDvtj3iG3kymIxURrwBNmvPUTIpcWxLDDFjL1qSDgRrl/0O7EFoFx/YO1gZ
RXXFWSloXsACihmiT+OKSwlK6ve0SSdNNHKJLNVxhMRIBN5EcQnD6wvnDiWbLYpd+AdwjAbTdijR
ipgTHhDl9sEV4jMzOILDIIUh2WMv9IxzLm5JWpgVCLYrSLXdLjSN56Kyr2mgb3T4ag1uu3x2UQ8n
IDPQMDZgUdGLYbX+DgJr5CQaFVvnYdlMEVyguBq7bbsrGkBRKyANmH/WxeSM7KsKjNuz+Bx5/WgT
0ckpIpqdOYhAmbE+LYYLdgiOi3NJ5KAMylIpNiTOS/YTw51c2Zef0jg7/bWz0A0gZCkz2iC23TDs
VS/U6vBKgVLJHTkZwEUPR3Mq0GYDZTXO49xcvjTmhcoyJ9l/33sfNUDhSV7hrpfwQ4uwosyiAsqf
olFSzkpFh9tqOd9gOtEIHJY3DwxJeqVmQHX5ULsyKdoPWFJOC+toPe5OP8rVlU/12tDGSL2QyP7q
WCHlfj0xvv+nnWEzFzoRYrwiuvHX1FhH3Z8UN+ifpBa5MUbON9djnS7zadBuQsn+c11ONzf1DMMU
T8uV6WYqYPwcZIMUldwmSx/u2nUQOrynSHL3izUz9mj2nZ5w92YsjttiaVb/JXgpwnnZ64MPOBBM
XyPVvE/O+nMzTsVrTzIVHin9lV6QBCQTiFrxzDTrBpfvHC6NPwuD8/eLd51xGYt1s2SMYSdTliqz
8n0av1sQvqNeJ+AOUdclmWr6Jo0pPJG0yNU03RECFeo8cLYu9CNmQ6Q+JixWVvalbZYY1pGbqHQ4
wMtG+taCTTfaxdlS7mgUzqoelXFyZgoVvnNzTI4UlCxWw4jWsAT5NbvoCep80Dhern6lisqSosOd
m/cqfFpYm0Z6Ey3pinkwAjYwkXE/M2ScTirWdWSuFaAUwfnCCLZe8pHc4ck+p07rPwNiTfdnc89y
UgnPDvTMhsP/3ydkRt97XK5JsvilcYMgsH4jSX4VIepAD8sSAnHFAd7Bz7x+r4zLQHJ0lS8T5SGC
5G8f8eSsQt2OUtTEkkQ1tMzZJR02fhm/fA4J7WYUKDZMMDhSY8Vmlhx6f0fS+0QR+mwNkfEM0Q5c
EQgAXm153AtzakouRPD8B1sXguXoumCNYPnT8oZBs/M9PGEBkYxyqZHzoNyTVFeySIygYNhqGTbR
Sbhz+uLN8Q6sMJyQV31xvVsbStIZ26JsPY5lPpCUjIW83uKr/7+ucuAzpvXT6oJqUNedv91Faaf6
j6ooxgwiwVM41XUJCr0XgZ5xGAsZ3DmH0mQPIZNWdxcVR+tiAuouQyxNeRQD0Vjtgvy0RpBoNl4U
3MTn/zV7NjNnysFJa90fjf3PC9yBPhNNxwQumE7gq0VRY/8rQbygHpCzsEBx2XkicXg/nGYjjY6k
ofkn6/mAA4hZPweDKylKdUvO7BiEXapo0l2C7PskLUy0WlIQIRppVeE/oWQd9OgZgLxCAksYHQtF
WFYu7Q3o+EayavKNIVKYMGw0dOlEkuBa20K4rBfog82Mjs/YrqTqCumcA1qr92efGuO/Rky23GJk
yi96M+hJN943u1ljF2Kcs02Tk3MI8uRbMQlLKtLfB+mbBmZ7v+3FgQAYnA4BOnsJF3MFjGe25ocd
dRoB5ZRy3Ww4/4jWQJzpju8K2/JSZK4Ud6ujNVuaBGukuwMPJv6xaD3YRwxGik+2v/2y+WUe1y+m
I/Gn15ZaUECsqv9QpJ/PTbbV0XGYHWUSBMqtVKEPSd1aXBI5gqwyu5+O06y20JvsRDknPcSRcM2c
aCcbd9//TsNZ9yfOyvjbuRIWFdkvz4bb9UfPaGvclIZR9NuRsjIS+PHeGdlEV3C52cTQ7xMg55kF
IAVdaKbSvf0tCARso1GSJdbexuRNzmtueVA5F3hJF4KSnGslEhcb+UQE6/Rs8aXvvtL0uC6LD8KZ
N/LEi2+n64NhVQ5GnTEWJVYRKHpG3WaWCQeqTBo82E0CJnSpDKtdziyhdAtrBVxNzWO2emm5E00p
Tr/d6VLT6T/jVa8UQik4HF9gHRZGZFSxpQxNfTRw2nant0/wmcqKTSSUJ8xT7oJGZvG0XPIkiKrA
wjkT05D+2iZlK8lgmTKsP08vRDk4qXc7cxtQK+pkCtkj1mmo6u638pK0+CF1HWRHyahEig1QlDMx
frwR7840ciRpVuex21u3hOmNXKZ+6zU2BwYZFaGY9sFMN7u5Wfvjg0AArguhmEzwmvuJ8yq1mWCK
/GYibGYHhy1jmSCNAwkglfYtfUQcCOO/2uYt0eDEmuSSwkLxYRlmZVY9Ff89KDI7rTLnQokQHsOY
GzMfPpK4GcIgvaOVHjvNbh8qhzW2jh6hc71BFG6M/o0PqVs+aQ81A1ccTMrb4SWiuUHU9cz8hREy
saxmScsPuqMnWsUO0bKC5IaeCTfX9rUE6XH7W0HYckiz7poewZaFw+W0CVDsHEmo8AlHFNYqgHJH
oTfs16oDigLIIbtWJM2x1lI7cGFGm1/vKxvj3q9y5xtRwFJF0vSJttziDmxchiMZRWvlVtt6xZPL
y0foxf6Tyzn+BQk3lWQFr1uyjkxhrKGKylBrWNgcZKUtWRTYVcBWZO6P4Tgpal22wF1bz52Qb4/g
4NnKQpAZ51r4hXJ2NI1F2zBoLyXwUCNcTdoGSLU4HmWra+W7a5zB3QqlbRCuzJzdXZO3TLhumsJ+
mCHj2lQ0cnODOqyrqLRCavPDmKw3Cd64JqPulvhQwmHZirjeJ0qRrRvrXfHj3f1XXemVjLkHPSAV
Rqim+4dwWUS6kgzMLNLURaYH7qrG6HnZhKSU7/4jSleIJbxrnPAeOTN8sq3L/gim5V/SVt3MsNm5
Xm2azIyhTktil8ZgObqUUpcMVs7KOYmF/Zgx8xEVvH9j62VA6jrlTYdU/ern2hkzStn0OJz3SXDR
LF4NvAR8bpPQbGnUunNVfs0ENPYyWs/uBwphw/5kLY77svRiNVgGy37lMMW7/jN5/MRgB5leKSHJ
D+ACe21EkLcKfBcYQe+8Y88r+kvQ054jzx/FKbUrgczAiwyaLKzbcxR9wtzFD2cehPuiA8Rt6GY2
K+r27BhSAl5S7U9PLoC0M6i2qW2BoE0F6GGALUz51w9gLqJv5mcldt09QarMZSCHLWlnsup7vQxZ
KGf0JsROmDYjlW45FvsOIN4crW9Ncngw9slXCS2Sf4M8E+DiXCuHYSzJM2LptIBJphmXjErL8ay6
Vn+7PKX5kvTYLFZKzpmpfLcbFchJuvkGwpbVk9U3c1ymd6q3HTGOkPItkVxuYMIDFMISdSCY4b52
x4BdAo04jhs96g/0j8owX4VhGFdpH4pW94Z3SvREuo6N5JDvnkG4YxhT/16lXxbCxK+Y7ZO/rHvT
ixC//93Zef+2/I0LdOwxpNna9EtM/ZoAn5UGtw3gry0QAim4zbYh0zDdggeUoHGFdTu/J2+VFH3x
WC6sKO+W6UMBDImbeY3bg7WOJr6aIQKGRFlmOMTJKScHX8R2OMZa/Ax50P+u0yNYIMI9HGOBTSGh
/g6Q3axVZnpVIW4jHVahMaWJ+ualkfjiw8T9RB/nYRhytFv8rbhWGAkSRanWwgp4n0f59IaR83w/
AWs6JcMOKjamjv/aP93TemEeltU0km/vb34CLOQz6thDrVG+hR6yv6uU7KljFNHITnaBpl/iHySY
DnU+zkbj/U8/qdcjWwb8YFHLC77UHd7LhUVfN5D0tusNw6jTayBO5G3cnn5VL5+z/tOKBD0C8ES7
tCBjA80wApNaZSf2yeNkt9CTGxH8MpMopPeijvM0gtldiLW7YmS4ZmF1humDX7xZ8CIUeRpuMFdx
ZElS4nrLWVkd8AZ5iqY0X9FDQC/9FCN6O909WT01y+BmTuzW1yOW1CAr/kMVMRTw5aYNrGsq7Z9R
BMrGGPuRdEYi5WSatOj7EjhJEjpBdRxgVeDLfNOrbGjWe+2le64nzDJCR/0BJT1BS7nR+wkvW2z5
aiG3yXJJ4YByjxBAZ1PiWfjGuEjEtzRVt9zSz94gGe6+oGQh8uECvKnWgWGXg8OOysvGoa3ke/Wr
GxW5pjgVDMFFaE/zsBUFyCymUkXW+yoHzevWY4yYzHx0IdQ+7px5Yyrd/L0Y2Fq/urZ8UAW49Y3y
ht6Yw2v4LKeIvuwJwV4ovjyJO8cVpfJy0a7wOrO3wF1rPJ89aZcgv0SNLUqSjf2RxazWfuo6xBIV
adRYmaW/TcXtPXL+oJxAdvoXWFwyVEEL8wU3T+2k6ctfPeUu6mZjjI6iydQGJ8Fv5XvSQBZxS8ma
PUrwBUJ2UCT5eHJthgwUdRhKL7TtiWhMBQhTXddrYBwkZvSOmqtYWbJ6H9WtpkZSoy5VJzwbMsdh
e7jZB1b9tdth8FBgIal9GyJu2jWRDfBkWtktVoU1KQDcTJczX2g/RKMqCHgXKBBrdKCV95UubVis
+u+H0+UAsTXI2/HvY3LQBlk0/s8MMJlg7acx2wZPjGEAX5cOehnIFw1KE7ezELazPqkfZwYTD90F
oxss7pPpfqgRC5ZdofGkf+MSY7AOSowFnvSVhmovMPDhOI0GBrTYfhhBLA8bf0sz2Xbl2/nIe1j9
jSFexcpjhmqKjgFGJs81j6/VkaU1KMEAQqmgWnZueZUrXj38bR1GjOy1LMcCo7qZzrAX4trEizpM
tQdqpojePDHwvlurCgI7dKKqhCTX5eB1u2OBz7ibRVEqpCFWxfGjgy7J/4AG+c9d1QXM1F+p/jwL
CgtMhemNWN9M9oX2fBOM5ykC9tcbVudEq/OsU+6vmyN02blECeIBbE947gk7TKvSkb91DtO9lw3b
ONNusAtFSWgYzVv2u5n3lPJoxIKqHjpprEwrxCH7fAQTgkY0iMcFGYuf0Q98iNOMP+/SFG+kvCTD
REbda7Fjv9mtAOETSx2tQ+VywagrBRLaqMYITYfkG3RoPhQmCUnYb2lREp/0atJIhFQ/7nFXdiEz
t+xLnLgW/aLvzdZRfiq84GtjhpdSV6wNapBItURH/73c47PrQf/QIgk2kfW27LMhNjocbArE2EkY
K+fDqhJkUk2Ti/Qz+8lhUZXWLuo1Ixuy+Mye0ZhBZqpYhFOP0BIVJ14AYhwT2XWWNlMBwDoBF4lc
FrOfFcQuS+tWRweR77Ni0h2yOT3UGkK+HtRpaQU51UW1BIp7eyEeCfJT4kZizftvIDW0pc9duqbx
vEpF9BTkhLfpICypykIW1J7KC9goDH01l/nj+2PZ4up7Va4VtlLCs6heMt5Ss2LpqawBMIawnuq4
zuMCwNmeEcBsfRZawYvgOjKEEXHikYoEzlka3yzNrPdEu/Tcqz/MvLr69N/Tym+DbgypnNMqxglF
qlx6rFjiC+x7YNQEqDgl2px923NvLYHSZb65WRlEGmoIf6Pv9rcGEYdetiQ7ida39Y7z5bmmj9Sj
L3u3b3HmCJEnAF/5SCSx5gd6DlilKXv2PkMZ31hB49lV5EXHTiWO1pM1FSa3YTZ4BlpZHqCCwpQB
2PUy4fs22OyqZhceuKvXdHuRA2Uy8+W7CrlhexVWwfe5ZmDcZv15kRlfiBR3Q5f/QXWo8haJzMdQ
hSt1ed+keC9VuwFHxg6loMGNr8TRpSwiYd6jfBqZUkT2soISv0oEacEm1dCwoctYEFLZBlI5gXtV
vU8YEn52AeMxEJYYsAMMdkde04FkLYxNKngqEQ4HAeEYOxQFY1AE0aECF9nwsKB4CMn5DffehXnV
TdNjfuxzse+NNsAXPNODxC5unnGBMbYC9GC0em279WoPlo0DjbArL58kuzOSi2Lf8qwffyRHyanY
aWJOW4xQ8INcuzZKKqWJEZ7IL46tWIZtfXMyqhQhbr6+g+O68KfHr/YmllTAbG3z0qPoJQ7B1kFe
Y9jhrVW1coJt8uh7GQMb3aEmbNm5H9S0qBVGfjAyi6kCKwbIyiX5dNwUzltvN2wC3llLebr6kBRY
Xq3f6hULJE9ZkvVNObBCZiBa39KkhRNV46c6fHCK0zUjBKk372GpsW7S0w49Cs4IbFJz5OJAHmvB
PVVZHkPvHOvck+YBB41F9UcK4s6xazNPD+z+YwFCVKP4/JLjEB41RXWiZKlA7ikl7NWTSkdA72IR
5j3/6Ta0TKaBNSo4Y85y+hVIsS3HkuA6+9PBmzxyACBQ9jo62geORHhcgHLc2bFVm3ouPlhSIz2i
Fb8Nb4bg3UOqAF/f21isLqgm6b5w5fjxMP5kdPQbyblaBEKUOiGftznnJWbkL6ihyCsoa2FoT3F+
GMLoopkrO5vYrEqkB4Hmk/A7xxhtO4jbiLNHQk154GjUytLhIN0Z42FppEdJ7gjJ+sV6qUlpQKqu
5iv5ZrHHn0WoKSyw3Pcvu8PByDfbbI6imaPgVCdYiTU3PPoAo/Vf5/x1KC4GCp8LRZD9NO6DMebp
idQgtuiYVULrXKBfB4pBHmSxyRY4SGEQ7nDLFsbE1sT/DqVMPHWZljIEM6XPdTRt9IlgVtdApBOL
2raZytERi3cRWVnE/9eNoABDp9E/FygEAoMm4qYq8FAne2eZWXifXv8dZa1HVDpcFaOe9A9aVRyu
0WslMjMdbXFffELMzyoULfpJSdVSQr3Oi1gicdMDc7TmCbFrkjz93WjW2BIQq6s2WObl71WXq8Fq
nTg9UzBmk4LBhv+NI3OKPeyVpg0KtLy3WzhDrdfjRTmj49qhM9bcBAY6/OQml5xS9PsVAHztU5bQ
d6lxY5NEIy+CjKD29wj/gCuIZa5nFactucC4+7cDlOUKbp5LVUISt6nUB7Kg9hbUzbRGdwm6ubWs
bhraKx50nx9r0kabeqgvlzvx+8er76L86rTG3C7fI7A5NtKTjFuGvRkn9nqL7PiV0dZs7MftY7rl
zOoDuE1XcnQDCr1DbmAy3LLSGtaRN7xieKJQBblpaBRSQ61QTV4awhV1y9rlv8smBTtFqQqf8MK/
ZPPLBoHFta6xvuNceEOnCqqRc4TM13KXk1tS2Y0fwj7+b01rg9wFN1g5hpD9jWZNcjWEhGk+Rzqs
nq+7bfpy/nG5mEEfNg3Sis9egUN+hPlaLe9D/90kaRHQFGNd1IptiivIhTHECpmziGVGAKhmP8DN
UaEJtwFio1Q4CLqensBw5Ji5Vh3krWQWGdL+Z5CtzrxdG8wvQSBge3FIabOmHtK6sVgytgb/2e8u
UAS54JA2sair0b+8L3Q3uAoJPd3QGXXARM1KzT5DFXzTnaktw8ca2kx50+F7/WSosk8bxltJPXDi
AqiCnJednMbpXx6J3Pcl8dxiCI5iiduuCIaDQ7dL3Pko2Ax/wfY4GSFYif3IIh/+P2tHfeejG2PX
Zmk7AJTMycgqD6KG+9Vy/Ip1IhWo5ByZFBmrS+KHYuLOHkhoOlU6hQ+hzKz1V0Qr0/5A+JwdsF9u
Cqh/2Dg/hywBGHHWGE3bFfEZ+mPa7BCi7IZRuVg0LEBNz3tbfmsY29iOUaUOBNvic5O9D0F6SzkP
4QeyT9SVWTAYyYXq4WvYyogZfJ7/yJE02vlqDCceqTSzdFD+hRBSEFfIzoQrJmF1YOC7VrPrP/S6
l2xZ13jysNtGQvuxPn/Imwb7LPPo/Q4KE/Q868psdg6h30YIw9IVUwUFoKOyZiypNoAukeOyqMXN
Dk8qU1GsnGemeA/mOnEmoO1c/kKlvyZIkk4lmtfhuvEeboZ06fi8W1M2jtAwAekHVmqnwWvcTfl/
zjKVDRu2Zj2U2dUnYmuHX230ROv0uZTe/paflfFWv2oKqwhUqB/uC0WkLkbFOJ/RdchYoRZ6u2es
X3YH56pgzDX+JWjvvloL5MeZHciYwGxPKG9R7viMtGBVli4H6GFreVhkVly9qgMoJ7Aomu9x7isz
croJoaognR3NNNAMS/r1FTanQVgTeDQ1DFhOB6JQOfihXO5H/nhIX5+xDefG7QCYq76PWoIWUHRG
kCGmr4B1fGsBLUOlThN8Vf1xNfHOW76xlXoEp1ky0dgtVSA2erWDwLELBLPNutgwFqw5pK1oKxVf
Qo3eDVqIyW23ze8jrG4z0oI2dkGoiZUBkjxebgsIyAc4Mb50C3VgutHLnZhOEtxmpdEihLAb3kS+
PwDBQ4J1mBV/Jf8wsJsQ3Ob9r25/CrP+yydN9NfLgxYt9LuEVXXenWX87EL/7A7iO0dcOGeaMYO4
xXpD3jq26vryLKuYeV/eIqj8o5rH+DTdv8TK7k7SW4MOHK0q62Bdr+Lxnpwutcq2dJCtaAC0vcFz
cXoLJjVRNgLt4S+GkR+SFe1u5EbRX4rUOb1gcd5IiD/1pn5Bss1Sageu7sfC0fOf2ra+DiFWOK4y
zOaSP9bpcgbE/WR2wR0YEM5RfwAw/n6tRKMMhC8uM0Jtq5LjoVEdVh+CaPpVwTiYMDgkivCbRndU
+/X1oPU9bsZF59X5ZghJkylNHrSEie8wnz1yS9OGDjEIE9WT4C4v0BonHZBcS82RnFl8e2yxmQml
vxsaXPzW8QnqaYI4wgYvZYtKPOrCzomU+umAoPXKPNdGVfMOuDRRhfBm7j4wx8vlegDnN+EHedfq
kOJ2PP6/73cn0nVJetSOrSbBp/MxdwFv/JDGcvXlE8IS9eLvOdqD8tQvU0FixBpHqo7OWvcuGqA0
iP61JSktzr/th9TjqkOCfp8AIrSkVD0Ci1HiKt5/ZtGvJZZgGvB9Vl3p1+YpV8Ja/szkWgqKhst3
OC2Jsgf/dRLRmMhdyS1qW2Q0vXK6jybN3s8Na5aO8GeZil0DAjVSQUsNBJZu7SIJs0genrFita1E
Y8yiSuGOEXge5T7po0qzTSBzxwKpMvxRE4PIRvPyG31wZ/4AhXLRoxdUlxQszF/cosexlvjXOal0
s4OXudNja2PHYWg9RJszOnoDvtQc6jwOR17xFUf07ba4PoLLZf6ThqLMPLsqq0DVj5TeeTqgZptA
B9RZxow78Rho6HDs5lISz1JBNRW8ZeVljZgzJKdXIYJus6Ec6kyMBEfYbAg0qQK2fi8e4HaDPWmq
xuO2KigDR6vysgEUlXCIMEKRSjj/jHv9DzhQiyePUN2kBhgoiaqSgfcnv2JtEC16nTkTSkZusugP
8XVZF5pDhp4DBKaXDU75pq/x4HOWAV97Dsn/dCRl9vou2kWsOw7YBOp2faw/jxUWZe6/2oH+OIOr
hjJ+l3gEzFKWKx2Vozilzw4EvNJDa+nE0sv3xEy5TTKEjo7M2xaslgyt92wERFWRu3ToLRp/jw3Z
k5oeZFlg7t27UpOrjfas0jUhH5nXlqYt7Om5SDT6uKoSunRW5docFw0qJhYT3h1o6wCuiwgzkavw
95WrU7EjUshksJ1Ie9+nkDDFkELxjKgD7wDR2ggYkR3h84ca5zqeKj7F7eBKBSAzzy7gXA1ECxXe
gkgWJ90yKZl6CHcvvhhV6an599Gnb73sNBPIyrGaSbDJvOZWbKWAj5d+jdHgVMXzJRhZBrSfG835
jHUO3B2a3PRIqYisaexnvFJbNYfvbQ5hctoQzJ18GtHqKfPw3NLYxuWYTlFUCwVmYi9YfMFHxROB
cCtNwK787aBWGfO25NucKyaEbocaCterSM08NnWnCMiY3nvGJhNg+wcrFR+xJ8Srla3UU2rOfIN3
5kvmav4r5xcW8z9kTkegwiH3aPleMZ10i1e+abiQIwmEWmZxtLbu8vBrPPjQJvrqUswwLqnA3L1Q
fNH1kgMvM48idoAxX3IHgQe2dM1D1kFgVMQSTt4kWg5VwHJjIro+ui/KOlsssPY3EmPlDe1BNjyP
bRFFlnFKVwnDYFPcaXUGsszfcU1/nrAntsuwVWlBDjTh/+rL6IKYw/dE+pDigbf7LwZvlwvE/Q8N
PCYqPO2qmGR6qzeUgVme2rZlVZMjAJIwgCI85vOxwY42kjZE1taID9UEfjfTwewIAgvvuNDzBWEo
LyybDUHKYh3/QGfWkZYv1i5X63rzir1m0d0tnVnBzjJ3TBJcfD6teDg1icK9gc0qSkt3FIjnb7hB
Hy7I7OvUW3nD2shAy7zsXsUB71fWSscdGt4GxRt8IbmOol8uTZsvjkh8ATZi5Kpr4wJHViY0Vyrk
LRl/rgAFoGMCnzTn9wfL8AZ8X+oBdlUVIff/U8zFjc+Xr/ADWBsCqCuafbg7nJq8lew7DJKzXf4a
tl2f4qa0dkvo28csJ8uXtNJznGQMr63eU2pocArC2Jm+fIdTg5ukwDFSVTNhHnbVNEYpJERuZijj
8I/3pbaMQp8gsvweJnwmxuaVa5HxFIAEW7DpFf6VIS+UM0wS5bHFe87lzuRq+Nv84EuZ9Cf3mSlR
dvH0lqv1QVrkiEHlt4FlM0/nY+R8Jk61NqLIPd4spduQFnLBWbxwfhiZJoWKAR6020gNrKqLMkWK
boe3ykTrsQWoGQ0nnsJH3Jg6iLYonP8mXDzn5JbekABqLyLsvgrcOpzoAhIUXdbIfAQjFctjYokL
d/Ghf0laqFI9gbTpPW4affE2rDYU85WuwcXmK4X6ApIkrK9+KKCLLsc0gc0TL+eJdvomE+DyZOPo
GqBYKcyzT37QNq+f/GQ3S3Mv+VjbzLlW5MIyyNQlTCPth5wYSIH6vEW5Fc34hrwNfPSLozxFkLky
PnWNrPetlKuOnRbWIqJ11GE7MqwUlZmJ6oFu6fCYW2bd6ETe4og/0lpProVlDUYaIELd0NHhaKwB
0DppleJakmiPyRNYvNSZ75jnVs8auAQzgUhKWXYgE42IPwI83PcqPxtNSFf6nE3ppEE9EEym2UM1
vciSQc6TJQDWHKT4XJliydcvvys1XU5mM39gZj4MqthF7IARBtZxjVI0yxqF5vN8/m4fmqmheYyg
Ek6gcV1UJ8is+N1QS6GPc4PlzskmS5DTzk0pB5tUYF86MpUec9J/okIIeaotwrMDSLWXqgVH1VhA
xotaBnhy61tn10rjOg7kGF1x9PwfppSun8OuRGkJLI7oteXLd90yH0Lduz25sGRVqi3poePwFbOX
LYjxNeAX7BfOAPi5BbLGPi6+8bhS9+uJPlVPf87tUypKd62GU0wpiXYWIXRDPbcK0jHDKQloqDcM
XfkK9OCzF8sWMjVIBGxuzWvBdQ4tzDgFO+6Zqf5ef8YaRYbRYKfOiTILJg/X3cKvbBT4Q6tLdqAl
0BjoJY+RRjs6cSTlXLHuLqrPL5IGqejF2oqr5Bs/hvrLWU8TyPLN+tSLTrYU4SIiekISyk9p2r9W
+Sro/qHFy3V/ZEM4VEvybr90Z2ceaXB/CaC5zV2LgAfO8//62XWNP/hIUVzb2OfJeRnZ3xC+Dvsn
0DLLA7aN0Z/FRBnDfUxwOWCwKvg6cu+UZAwrnr9Ctx739xn5Cp7G9sLJVuQ15kqCGcVzK/axIi9X
U3FL4MFJqbldu+ioKWZ0r+L3fwQx91t9P6n/t3wWRgqgKYRvRn1PMmvIMYXI7HMMzWfOu01Ji4xd
x/st7wnQeenwgpQ2YA4VYOFB8r6hh+rosB+De9CgZn0c3jcbSI4nj2ybgZLrFT/IXEBe4f/RBnaZ
Q+tGzFaNcbBzEnxVNOf8jxOma/Um1+l083vC60jy7q0JJiwQC91AKBuwId7y08CCEICAZHNNcl/z
8ZL7kJwdfCkybst+pjRlBoIQygi0EGN+UsDwir5z5DJ7C+ADo/D9xla11F5i2e1PP1wHjNrF2if0
owfjLqqPjI6F/hqpM61obhUpdXYXKn9mQFgBIBrN6KYPXz9CPZHbAddP52tKj1L/jc9Cb6exXuWq
Vo1+IB8XX32i/ihB3aBh6Lqx/nvpYrDeaK4Q26nAlq4yFAwiT5gS6WjSG8wUifPWRyD52If38Ld/
ktXBJYdGS5m+gzZ9ec0PviSTuul0fWjZHiwlbIZRb6tuf3jX2nGLmhW+aqbmvUgyO88Ic06IHBaI
lBUAowAoNm2zEtIIsj4PZtUwKv5zk47RFaJo6lxRaPgGk9WGSTnxfaCYj0fMEixXOmqNpaq3nnn1
/OTReawLb8dLCmagDWhH2ydScDi4sjJblzMK7q9VtP1klzIm2j2NWpOnUTegYI4jzGnHQMhe79Hd
uVIBrIUxiPLGOWLQ/d64nqCacJW293z959BtP1ipMOyXzm9HT2q251U/feJU2fGogY7fUkDzC3MQ
sBxoGP9xTVsoNS1SEti3IwEnjuL+3iipCS5h3I2xtyTsiXqEfHA0b8+/F0vyo5o5BAodyWwRFbb7
nKUzEekxY8kwMjm31BLT1u3HyLzJUpnDiAwQQ2M4uLYzqQH5zNq97Kg7k0amB+/yerN+BRiggbPm
2XG8hU+1qVFX59QXox7M7YTYIXU8c5ISHPN3MbvscjU6ojGacz85J51KW9WFaUM3jG+ZTMPAIX1z
EEjB1BJf7jTokIWQw6BVXRUhaWqfnEo3T2TbDFviy2h21GSsVApTfVWP4FGd2Ebzr6lXwbrWyt/V
wmb8SXXgv+iKWpsJzhPS3mupW27HR6sm9aZadcQ3qTBUG1HY2aFLiXR154CVxJa5vW6VjTtZwKPa
j2f1XcE+cmKtWpEJzm+EdeKq7gKKRG2g+sn/za2KdFPZn6ITpwv1fJcmD2ZcVMn9+arGisuRST6i
69Loa1ybbm1XJnvkgV1YpzfDAgFkOIAk3xQhkX+vd5ndEZ4JUuyDzwWkTuP+u6ISI//CoNjw4iL2
K33JKKkf9ssKhvvGkGdAf+c9bKLqNjrz0Du0Czcu8ulegr0OFLV7rNU4i/9okFqHBzn3D77Z7U7E
alnvUNS1Migqnb+HI9aVE7EeX5G74LkjN/gcCmTX9Wlz3tibxjSQOvdZut9hJsao5cYoWYVZmIA4
t3Mk73VCF7AwKL441lVvobB4sZApdhH87ZOBNw6ltSpaaDMA/7tXI0pHZISffUUuNLX8vol9BHf5
zLH+7nGTT/B4ZrDJIGlXrXecqvIxU16FImTPMwhG4guJRCKQFc4FpJjneN25zALuLpB7c5XOLFXW
GsRBSHe8BzZtU8dvniGdIY26uar5ovXqOPv0GpArCJAXzgzUDD6rBJuGrdzwD0qGDiCGuLatV6z9
icDkoRKfC591w78dhzS6ANWgL0fknj+ayr1o1jUQjshb+R9xEgK8QzYMCC4TTDIHT/1uGwzzDNox
bmHiywsmw4mkuPP6HWogBsmOIWG/ue4QzntmZblWFY29ochQzY74ZS9KW9vGF4s1e7MMvly1YXPb
RDPdh3EoprtZOUio7Hw+0ZSuPSvSGJJxq2y7ZnLiYYLNdHIVLDeSPr0+13wrtwmsd66Azqlk0T70
qgr2SGYeR7jJg0YZYc2GCf2kjHo7j+8IuDRtbFJFg8s3RybXzrfFny8JkYdUPY8mdnBVlI4Zyw6q
a3Eg0rcZHIgV/NEk85VhTj+qyg7y6hwCAqvDUWTvQJeGfEXp2+pU0Wwo7uk61f6digzw9NOyE/rv
EquNnhnlb9hmnFM+dd5TPIfGbtGB0EmGQj6SXK5VD7xaejqVFc0CHN/uYN6wtV2WJE2uBPCK729Z
R6y++Z0hPd307LQe1RmHpge6/Vltg+WBICplXmyS/K1tq03sEDRdI0h/OMsYUx3xMyzXxnSfJQEm
yxUElubMecADJK+beX0mpoEuh3nNLto4HhjW/g9Lni6dt4dI0eow1eovJW+pl/B8OZ8G02Pad4qq
TUAbiKOtbPghVO4toTE/HPtOlslpDxEApHifnD+jZ+pFqaRdt1ucCUZobhLBwD090pYRC2nxVh75
+IhE4JLF5mQqg9PaRxXCwa9f9rFNOD9QGoWN8BeB/yt3g9khXHQ6wfJpJNWpHMo6CbzO+kpAKfDe
MUNAbukyVBBmU1tUzq/N+J4ak6bUsDYkZaxgAT/OajqH8KiBYZ6DWFVFxo6sRCOLhBV92Jr6Btz3
tFhd67EotGu1fY0ie+A7PtU0mRnRpu4LtCPE7d2VAByBloVthwIZrpx9DptRiafQ2u/rl87vmNcX
vAjzxvSF4RwISeNBaUHTRiveQYTGPqTEuGxUHSxxRtdKtUmoYjjMR3rQxWpEL0jua7Cbte5N2azp
/pHcNVOXU5r8XKbUw+GHl6v4S80NbiwbEQ/RC6GutIX5VkYsSqS4r3GCkAFAespZdDGWWNiGGwSz
RYcH+iOXluJJbXQN+Md9N+jWcpF3GFXv7zYdp7Kp9hjaU4CxXthgq+alkiy1lyfVfoCHJhMZuKAT
B5rZwpzt1gDT6VRcVytIyyyCd1nCcvt/gMCrMXIHUkrFaZyvl27OkCw7guL4jPc8oUB+E+Rxo7iX
ackPxUc90j16hAKXlF7+5tCS1KX7EADFUaeD5SbkC6/576qTq4hXzJxATp7Cchad8g3MnK/+q39l
ApnNU/osW/HjMhBLU3pt2FWw+Yc6QIaXLQieurm3VPYOp1uMTie7QTmgvnXswZyQo9leUbpKNPF/
DSgpw7yCFxcEL0Xc8fN2bC/lb5mZfY/b+IEE+ppCdzhcFjMyknUWS/vMqdabimooZPoaMqgmJK/j
b4gs64nsGdLa1/or3bPZHO8/72E9hlttnhkLVYG4Tl/6V0P5f7RFJJZqCq9vczwp/YZEAxCgDBUV
1X4M9aQsSXzV9UZWdxlEjch8WV162RvfEravhcCxeOa9gaAfUvWL/U/NfhUkW15MLXCBbKeXtoyI
NhPVz/Q6pVfx3DQcdxP6s51W72FbRRWiCyQOx5azrLTTVQe9totiZsPs2FT9iAaos9Ss9rAy4HE2
mkbRwvhHHP3RxPRofcBSKxLHLjOjvDbRpMUJfv259+d34VnmSava3zwlASxaPF1MGesVWl+6iDfb
F+1UslQREQ1RhfDXjzSC4chR4PQMhkTSp8WJ1dtjJxxK61WBIFAzstlv96FK5Vo5fump0+eSOMUV
2BRa1qJ7aELUADL7F0sC9vkzpUX7S2pGQb4li16vLQkR8UEGFBlMMbArtDyRuVLRk+Mn4a2dBENt
RL4wEtAGvMGLWEQ+eiumB6ftcGlkGYhUdAlGcjHY8MXK+NZqNbC5AAv91qTLXHpxOWQ5Hu0uOgKE
sYDtT/3nnJ+SQzxxnwyHvSjukLlRQC/st9lLK46VvGGj7Bfhu7LaP0aK+S9Q+2RrcL8DIgjUsUtA
JKthJsK+Ke8FEaylSjDDDfMAU4MSphQYqjmqiqHeHlRwF4DiGGaKJgfzOz2WOHctGLArRCO3oOjH
zYR2L+76NAHfKIjgOodvrKFyyRBcbftn44Fm1t3o7p3JOY4+Za3sv3f9JAOMFANEXtHVeUPdhTjM
fi6dMPIaTZOGih1qTL7kh41xQ6BlC3/OdnhKuwQR9+5/yglJhfZmbeC1N2sccq1ROwxAvdRicvrX
zrQzV5yeoR1RRP2cyqXtvdm6UHurgiAm0QwLzv7z0D6JJz5w9J7GJBMxTE/fwEx1JTol3VP083Vg
PkFHPfhbWme13YUv1115sRL9T37TnPvgnsYPCQmMKDd3ekaLzZWAMRVP8b9ulI+SAEixW3j6ErC2
cTV0tF78LeHPl85CfaEsD41dLkrDyDxmQCJRCCXEnfaII0/Z6f++7AICP0Cnz7tRWx+HEOyOtJO/
mKI68pTTd9d3HMaOIeB5wp88yeQSnGiyIs42jq81t3/oiazWsRpu4cjqLDWsuPTL2bRAtkqwPDEh
vgufnRicywZs7x6W4RNQDDAJ9JReFFRrGSHDjQXZ1Kd+hEU+7KUVvF/8m67MB6k5LXB1tCpEFwud
ylepttHLoh0WFOqmXiATvWqHhxWfSK0Hgnl6eM3GAqDx0YjBR9/y6LIJsUy78qYElLfvX0w0/4aM
zn/iysu7V7fduDPiLWcvXrqhkIDK60lQbykIM6BR4s2mvv43NyP6P24PfO7P6xwpCsOr9MuiQDiM
NvTFqxvSqURJPpgKAD3jq0vw7XUv2odG+tr172AO+0JrDqJTOlf6ZsjNfPuPOrAcvfYE0xyp0Knw
CMgq1BStwyiuu7OujQvr1OZ/9fZOUqaDiMAwPjVNWln0DPcXDopboo3z+aYO7zoENVZt8IF0Zdp9
YIzVGX9lLKMCsS5go/H3wQzzLhchnSAWy4VwZltKrwqXlhpF1jrQSCzSsefMdBbNA866KYzX6ODq
XFFMnYDhNJyx7NoVIDbY1j4/PsjUY6Qwze9PZjCVGEDYex9+B51QOqb0+4SPLX8nAZgvUlQyGx35
rPS2hHd2YK7ZrhTbuSLxEJP85VhllluhxuCpciYNV0uwjssf+kSi+8GrmlCmVniGOeXx0ddMBvWc
39kBDitZs6WZPjQ68aJhuct7cLNDzYvZ8o5pu0biioRZr7NSKKzYrA4Ot8DbSWqRsf020pIADMGE
ZR+b1KSenV1pD/oB+gpXI5m7JID/VmEQAwPuCB3qm/7yYqjBWBud4vxojUXn7gJWlNqAIqdZZj+b
PCgVd2TT5L7NpYIi/Bk+HJECUYIA2D62fLhHgM7nBr4vNYOsAMVXVLGe8sfjMBkdc9qdY9B7FZ0s
Yy14wp8xkRKWNnMb11bM2xAwPHXFFV8ru6QUx31xD7SKhcABjHp9cmChRSCdcLO2ygJPbgeEap8z
NxCP1ozw1pTQUfR9lNYQM+hLAybU7v0k1iV8wEOINyN9Vk6E4PcVvN2flDTldQJFDTxMEt80IsfN
3ZDcyimWqlZ/dElXBUJ4HQGmkYQEQDP52/gRTw5F0WRUTkMaSDJMl7T7SvvDAcnsLcDIo8e175sx
ckCatNZ4pqDQJcKoQpjD0utOHDQHGrz5J8YmqYyLg23aGrEXq/cwylw5dEu+udRKxaCyeezo0pXF
dxqchv2eWsO2fqDwd6LiLYOB+Yj7x3x59ptqq9gx7EMaUdxQ9LvVjXrp7f8wTNVOCGU2UiYSOYwv
j2fRHZk/yh+xHcNZv8xS53mh0P4jomJGnTtancByxZndfnDLuuwH0fBWco50Y41enP+RpNlvz+F2
LDzxf0liobOZ5qH6AogRow0nzkme/ldh0OsbnkngC5HeXpZ/Y3MlZhWMKHaf9anOYwcf7Umu5GSP
INeFG5hyPBj9i28KbPn+s1oVVC87YvTVA6LN2Rtjd/EDHfBfuhh9bgCtIxCGkWG+5MlcBORrNSrf
AA/bKrW2jmTkUwlpczSlkjhcG3tC+fjtUw8NL7AzCz/+Zcs16iUv0U0I1FGqoL30wXgzujDoA2C/
2dvSTCymWjxFUV1TtU1nnhZcbn9UYmnoeSLSskyI29gpn94Gqz78Lm9OkBWrWrFiWAoszp/0mJUI
6VNTez929hcbruJ6TjTMvaPlca7tAkiOO7e5nk9H1cGcv+gsDjpxImXz+w7xODUFmJFpREzaO8sL
gfLRlZw1IO9UNFkb5M1BcZtRzNtMQJx690OEJ0NDiVgwhqxqjoGlTlrmEAr2yA1OABPdOVYbHXiW
lyc2mgRl0t6xyvmE3RDb2gaTku/X7x2NjsXXUVk19y5ol1jBpBxygfEiXWuBO9stdBYidQSckNSj
hV0jfZoJd9ST2ioNe4BLpV/Q/KzqcgObGqWX3Pdy2pZJaOODAvKFKUptUJs9Llrvoxl4ecPvvmt+
Bv3BNQHZfeIp4JfYvOxlpXuMQkgKOjCZPqtfIyDLcZxoR3iAP8t/JfcvlJUimJVe+D6XoaGA06dz
G1H2RTP6xKrOl5zioyUeLbAKA0UU4yg4fltyB4GXLZYR+19mIckk9hPtkvpWT5OZdCVXDV3MuVcZ
DaQiaKJMzZDq0jq9TvzusgABQjYrAoYfWutU0hREXMdGdrYZHWrNQFB9+IrbhfSTba2aJhOtyGUf
Ym9PerMTek0isZKdXa4dluiLYCZ/bvYgUdZxpnu5dIUy1e3dEDrMcBwI5KmupsIU4TaXGVNoj6DR
LdEkumDoe6vzHv2zIohzjHrwPbgsmmHJXZSSPPkKVrIFvr7BHGlcSQ00cEw06UWmSeO1KRBz/QeI
Px+NMmUehtKJOppmFXM0+zzQ0LAafcypxV2nug06C7BtsX1EsgUDfv/lqJLKmWZFfF+h3KlRG6Rh
Wv7xUGaSPBxHVR3Wh5qwhjAsSoyg3OuvSrfNSLc+AKPEIArvZaWVMTDIaWk+kZPRsQnzbR8mOkj4
55w2YVVnBFEcL2SPsKtazIu2ZC2y1WvSbMZonxwUytP4VjcsRcQCWXUS7KSHPjX5oXHf0Dol7KkR
Kwxbzn1yx6AfPB/EsquDtxq14tCZa4r+lLT9/NrApO0zfj1iJKukezX3uTEDr0IavghaJn4kT6kG
5eTrgZLif/mwROeMZum8iRVTKwkcV17jdF5VtDppmaztl9fTFbsJlujxWgU9I+B4HPNUiCDInscb
mHSjp0AHmahVGWrxPKvJJBl4MKJs0F34rnyCuTMu+jX24bPos9WGNLvrSKJVOlBFEz/bBtjfjB7q
E4ihdN1Em30IYPOzbT6vDCQpem9QWTxE9BpcCMoQ77PwzUM8pVrFEUn7kg0exaQfmMdz6hDnSslh
ScFweAcX63TN2tvgt+Z+X31opnZ9nRdc7Xra9x8THn2GxzwAMtHRpELtMvMZgcxGaf5B5O8Awkxc
CULobYEEfBgj/jVKHQwVOX6y7evC08hIKESGgt+QaWsddaegktZzyH+BzrTZQISXDoEE4PYsTxq8
67bB8ivGUhHcsZ4tm38a3mm9CKrFrEvivMkXsoEGPvyxIUwZY3bUrzF0XiHZ/j3/byFGgydvVSc/
nmJRoG8lh2EwU4dnrTFj6wW3HeEqGy2UWjjePxULhZp6wPnMraqTPCgye/jTB4YmMb9IXjhi60QN
OqqqugIZ/Fy/4huXtOOZ4qj60GNL06qid/ULEqj6T03DNlxpk2EBZs/M/drdD8DiCfFhcJXaZEWR
cDe6FuwnzT7PLeT9AQ5zuBww09KjeXhofn/thrdRCteyQinF4+o3bm7lSWOBYt1sRtJc14qU7Ml3
/rYXWNT3bL6cvB5m/gh+mtCtMdGzbPbgJNm+TS8MQ9B0rNJYnZriWkSLSrRyVXf0fqS1nmMCc/mR
3HBcWXhcGlILM7FBtIA+Dt5ATj9k+T/hvt5otOz2aL7wtDMhTCfmYkgKzZCDKQBYwC3l3WHakvbA
OZphawO417PkJ9QBDLe6bFO3DvInVXWMLiGxjJkN7SIOrfxF+X82LMn16HI2HDfHPfwdR+sd0BeH
riicBkzE+PSbQaIrKej+qwk/jhIQRr7wlbF5etJkGcKT0uvISzxii+weUVH4mFA5YQeQGZpdE2gC
InGu4psq8reEcjjn+hSlEIbSh5ltzddYSF26bpY6MDPvf30MeWSeNqyBmsBXkL2v/dg3PuqOIvno
qoxi6xi6W8E3orYevVWAjDT4aS4xt8ctMe9EJomnuv81R15wcqn2CliNyY/pGU4vX86imKcB5dGB
e38zLwDDjj4G8x0pZToZio+D3WzWz3cBmkzzjMAfCLJuI3SiWjMaDRzHY800rGzuC31uN3mLZIzg
GhGdwxWZtmdoadmRIVxOXSBOjRDUZXFX2yFpk363rgLzmEwZoOFejKQieBW7zvzgkNWoGgWiGbzt
sYZE9vGOk27dAtZi4+dM8+a8fIPE6LbStkH4Y/xPmyRNyotgoJiS9QYpdiSOyTBANw9HS86YPUaK
eR69KlgwCmtDTsnvvvlDGrqJmfUnO9crVrw+NvFft4NoCSDtA/b0U1U2r0AH/chLCu8ewvweb+Uj
bwgy2YijDfNnqSaQtxty36vC4OJQS22y4KJXOFMMC+nDuigyUdURf7JUjmgmJMGa/n2xbr0I7Kaw
xb4VpwlABGpyX8lQV2Hg1HlgqZmslyhQgXvlBi5tgaRaeQzIVhrM1vpbbnWNHHZXVGgOVgeOvvLw
qhHmQwcfxWM3wF1T/0oyovLxf8rBFcgLuNqcc4v1o0dcgEIDwhvmcOtjJlKYVx4yQPasvOasrFM3
bU17pOaByJ+6AyRDsZjQQAFcy7LyhZT4EQoi75wt1uzMHRcKEOBQIbXizi5iDgNScBTzWEGK8wbD
LSmINkX5RhP3i3fcsF9fgdu6BzPn8qWZ5GjifdC+j+hX4gthTM4o2EkmNU3MmQ+XNhRWang5zE2d
/Xxm+o8HQ70sMzZElAXAoj24y7qSDK/wLHNhKE0vsEmFX0Zs69W9u+fqTsQTJc6MNfQyB7fdkjRT
NBnaesILp2hwXFQHYUONCfNwTcM/Ue45ZVOZ6BWdxw4nI3U2oe6T+HuUr92Qj0X0hgLB4Qpmllb0
eYz/O7FKmBhNUT67dI0eQAQ//jZmi8XR7j7UBnqu9yrv8NivQy/zPRRC/phN2u3wkI7MUWbUI4OB
YIK61jI1U5ZvIlUpX8eJO3gMBAlTkt5loNsyThmWQA0KLtj8CvJwZ1iyF0pZ7I13vqVLH0JBo1xG
DiyKIUJmzkjMieOnnPofrdTMaMfJ4ydn0l/re6b9QIJTVvbgPS2ufv9eseDg3j4JEJhF+xG0Svej
uSDTSISx/W+gVCWV5XkSSAAR1qro4SQwE6CN5yco7OCaZsedInA9diVuhFsmJVZaV01p+gTz8h5I
YvTW6k/klqULUfI3SwQQfJVtN/b9qXUe1RvpSiEgHBvj5mkqRtUGTS1OygjbONe2I6CuMW8wdUXp
mFTS/OPYb8UYp/giEGxPecyqN2Z2K9F/b1ibncz8GACkbzHrQ3mggnYk0+FxSzDfkgoTeNjJfnu5
UnMmh7HIQnpWaIJq1MeKz2CYl6rxrPFbp/Z+AsRJ85UzLFv59x6rg4/rzrk+AUYkP0uIQrLBz/en
8swk637np2e0LlshMxQhfUgMQgcuoNpSGUgpKaACfdGPecD4guv2jW62TCzrTPBPb8+b1ezdu03x
Curfsri4J0nOnPFswIsh/EEIr4EwhxjRMchlvQavqXg8tL/J8PWYhYm5M0ntT6PQvq1owliURJbx
ezZD8mz99RXya7inL8r+SUwYx8DycRuIxe7p4mTsS9w1d0OedONRB7N7im1KucsTKfSmXoVdxkeo
kJS2M6ZY5ayeAaZLnI5JYkIFkbO6sKkqP0iXsQvOhscd+9P1IuRJciCHbnPxIWGLTcFcJayO4m8u
3nI3Mq3WoV+5aDrvL0qmU2w/r4Wn9vY2LVvXXzXQLMOHXfyh8MOjUQbTlSajswioIurbMQ1Q86AI
Lwv4Jke3IPhJj1XhxvrMxTo1YIpXUTIR3+fItQPPM1rAXN95sHI2q2ePpI96kkcuJNvQgUkluWAd
rMJAtAorG5a4EGSzZu0TKSiPSf/NtgMwY21sv1QI98hvqWQKJNgu4PIn38Vzn/WMUgupE4CtUQjU
3He2WKZIvhPZuEDuh6LKUk2caTeEmpB0Cb2LTwk2+OlpwMWVhSATmdTG2JB/xxz1x6OCMr2tdH00
pzVRgIFyJX3fLG+s8E66WNS/Gj9QXyrZxbw3oH7y3nuys7Avnys5vAJMxTyg9r2xnbckmnhVWGpF
GQnSlOOBVC/cTCDilT1jh7s8yxC5Rj972RPHolnpfpCid1Ojcpts/20DDxL7HfVMln1m/I7fm1Wl
258YB4VnyASBRFYlGbm5Vi3CCJ3l42QO1KnxqCHXuvJwmOJepYoNISuHqamSCQ7HUVlsINk4q34T
iJxFlaQ92C0LBMitgc75RwSkGhK1KpuTFo4cdRGZhYYWQQDymN3QOgUN/B64BUT5FOlmEvJ5PsEs
Lh1/E3uhuU6ZkXhKyd1k+I4oYsbDr4BAjrY08UhulA0lqM56oOW5/vNHz64jOT8V2LC45G/dT9HU
gBryGgkbXn+dNZJit6rygLli4hHHxjQCu18Z7PFsbAOZDI8Blt9uRMY+f8y4oAFgp3GlMd92K26B
6OUO/aOyQz5y9jSTI9LJKNNtJPefgdy2rDSuf5p0UNKBJqpW1oOxgRoJ9EN/9+64FNk+DVX8Q8Cl
Wq11OlfxRj5O6YGyCdnFYsqUc1lrdJpGMtQB0BsfwDPRZcXWRKA7tfhw2CGGFs7/k/5MY1MOOQ4I
wgLszFRni96WH3pGsgbe3iI4nl+6BMZHehUfpuozNi8nrGffTaMweVQh+6pj3Y7nlPi590sNb32J
G3aS7aXsDCqFygytov0LqysxoW5tGlcqWawBzfBMucP+AJPb+IYYX6OlEo90c9gQxRp8hGeEhEva
FxkmHJZDN26El9Jc+8W+9A8/ZpXcEnxiL/hwdr1ajvp1Ba7URLWmg6YBQpLGJeobOBjsrCirq5MM
zrxBtKOEbq4oW9rVrTv+3uHyCnk/TbMaXWJwNybP351W0eXCOLisjd3vwkFhR22OIAFTt++xCv6u
hw/IW+kSQcmcTyM8SIuy16/TWOlQHr0bilJ+FP1LC7RIiEGA9URT071TYe+3KTeiuSTQ0oA4LD9J
KrycQFH7A7Zi4Zjy2ScA0ptZFQEZK7CWHIcY3O1M31K8Sq6tnMGjLoNek5p15YYoBEEOb0qBLvcN
b8Unk+U+nTIgJJ0niC+WGiR484dmb2IpCKnS1Vo4Y3B6GyMwQgTooLYisYB0RksU1Ah8W/xEVRJo
16Zo25BvpdN8meNjOOsmbr/4LkHNkGLQ0QuFJ50E+lNUjF8xIOiyQluZfKPpYgwvEvfW3urZicak
eJZ5Hua7e0uhTgnexykTG6oIR1V/dzygDkIYUxUSSLpVmPT8iGtvW8AjV8M/Jafl9amofe0RdExP
hZgxQJXZgLsVkzJhPkfrp4ku7tFQK8wVtrqAS/OZChNuEIfdCm/5XwCrroH84Sz4vl35K3dBcZ/x
TJFaIDgqZQJRbzgeKKr8XLr1S41FxoNfus2DzBFHH9sHbvtRXxAil7rJfelwBnYjMtvNfBYKR22A
euMs127+ezi056xqq4HimQ1we2ZpcicanhqHStli6hQGyg9XmyNmI8p3eMa9vuiIODhx95oF0vqi
9tPoecXyS/OVtxwL0D81P5FpLUKX+hGivdR0sODXq8MFVBoIxtZNKTxLprsHm+vOmPnbideTN5/9
nA/wRx5O9r/6K0pWihnVWtGLuxbbVl/zug1amZ2aEbaGRILhvd8kDnswiBGI3blg7osrnbh5Um6R
CWQ1IE2paPz6YGg4J6/S6CXHJRbOIj95zJRueHBSw/zNZW1oFUfrBKszyb+35r4NJOh11/lNznK0
DTNLTQhkKKwGm1S8kJbYzs9kxFgh0NNzcp4cKOeT1eIQkZjQM3nn0b4+wIFgYSoE9GmHUGq5EeIE
4Urw3X/DPRP0s1bWPM2O/vGtQmnst5o5AOXP7ZZW75wXzMeJUUNkJ4Vr0Aw3v6SN6U1kjP59tzlV
aAmFbxnDJ00L4ACpIil6lS5O9EH8qR064A6CHwIMVm9cn0XI5MJPM2h/8sVtb34d11xcqwk2gI60
2wsblwwqxnkNHSqdZAEklwazIoHMWvKL4NlI+8BD+Hya7Ml5HUS77nKdw8dWx2ONkkU00FR/VUBG
VieV1tlgWu/A9UdJTnitovvAYNe10LwwhvacyZE3gFb0V2fsSMToZpwbTN7Qxvy6creb2z+wAdjD
FHIjkdofJPGrK5dkz+Nj6YKs9DFefGtQRMVeykQIdLTJq76yPGwhEbVyg7ixX4T/9pt3AaCk+2W2
pAIRkITLK//2A/lrl2qO9/hgckf/UitW+xrwb/tOJh7Q8ssq38v4enmpJ5qtKFYbWG6ZibIds6vy
BYKpzSN83RwkWzgp3Tn4qfGFK5jsDPaDtglJYf298d0GcrAMNH38URwV4wjuKGRa+qVc52KzT72e
CFK4DvttWAI1zf8ltLQSv4JryiA0ZgG9KqdXCZ4N1fJOBq7BK+gpy/rUYBvlhSztDpT4HSH+TgvJ
ZFcex4c1osk83B1Ignz0ZRL0D8MZrMS4zqm+NNrtsgOykOzy7AVgr9XgDuvCGJdXBpUbY5lsM6S9
qWoEMdmbmbqAWf1vHqg77mAXreMoggHdOYUyzxqdySCxrAqtuD0nH6alcy0m6ZwJyGThaJJsj+3E
okrJxO0mV/RiGi+cbHp5HFERQSNRhxFZhI7g6LYholRYwgboN7FU7KTBCyElxjIiC3B6O1iDki5H
29mf5DeHqJyercgGD7Q6NQGLKJjdLoFIRzRgXEAmCglw1df/pAkgFvbPCX1Q9CrA4DTgGmitYADx
j8+R68wjd8L4ovH18CAw/usVur7H9N6cZDZ6MIqgFoWo/G9C8twJuo9v2RZOgCsKOrIv0wWFQqwT
Qh80vBUyecZpO3yxdBIkRCXtEc0hpmk3geFj/O9LAIHCWp/rcv/BbLeFM+KRn4U4VRciR27Q8LOK
cZVSlNntcv6OeADa9ntXcYjEa8D8jOeYT7L9QpHLgssFgf57xizNw65e23vsTmZAaYOzuFsK/aKk
PWIzgEaqFTcuVy0+mhw+AiQZinhUvN8YWBCLYNqqOZ39HVhPyb9wHlkkaNp6Lr3xdhxMOkca+BJW
cEpKhZ02kbXVJKsEq5CognWtVedk9Wf8zUke5Sloka2opKa7LE/sYGl220Q2YAqrJAmtT9z+JKfE
o66vlHsnptMzBIHQBG5+D969rbt/CzLmQr6ldVotBMJoE+5JB3TtiEAGr8YZld3lMGE3Iu+DJxch
gRaBjqNF4zYE5wVmdEJ/HtyDlWaLZ49REu+jp9vxep+FIJTxLKRwJZUYKMR2CDlEGsNalZu9JsdW
BTCkXbyzYvoh/Rq/HYaS+NxYkx5NodgzSUtEtyqQWRq5e48Y3VUnu2IGsnPZ1cwEe/4NU8+zcJOr
qKQ7VeLxF1szctS79+9qxlPaUuIKD6kwG5T9SEHMw/CNNzo4i2hZmeoCEjS6vZ7wO3O2JQKW7t1a
vJ7Oebq4+H1kC+iMlxcSLO2o160rZ5KT7lIG2IQa2o7Qg76ke+1XQcXTX8bVA9ilb46LzY7zeLeS
vQAYXk2TcshuJ+8hOwDNMhdOIzLlDTQ6oaLvQHcCRwoHIyp/t20o8s2NrgEgDd2JagU4z490DeI4
QpXRo97x3E2pCelHvE3RhLWoMlhIG9o9/PqqGk827l7NCPgZewEflu88BYjJcWVc3aXWSKIiiNKu
0HcH0tMpcJRvvnRmf0XgZLtrriZ3jra2fBN+bWv/QrqNFw1ywXanY2yQFbsmIuugxUhjUIvG8H88
XqWkNrIcSk44ApprWrlxQyTcf1ScsJW37gRLLg/gjZDQotg+klJ8k2MiFIc1b5BwgdgEBuyRRkwf
0k8oxqNn2+CaKyK3t+PJsxhLDidy5fVkOjoNMuDfPG6outo4U38tOZJrPSWeEzjLEwdnmFRXkXgP
6VJhXn6oCZ6w//9BCJHk5vu8xTOtItZ3XHGMTF86cLAerSqeGrCalrCwiaF3i60Zoy6LTT7NIlG6
5LlHoQ3aslEfVk7Vq6ZNwU8VovgpkRtAw0ee2tP4bWXOGkhduHjmOcKffJ7Fww1yRkQdJRFNFlFu
BoDbQDgX0EKJ6yaQ4jgMEM5vU4QiF2g0wkQ0+TLioXKeEOpPxIdxQb1zM7LqdVxQBmdk6fW90QGa
aL3LmE7Tl22P5G3o64c0qOHYkuMJUy3K5T464HqUmhq/WNfb1cO1cAlNVyvaEN9QhbGfTjnqrb+e
jXu1L1cJfYhmfI2TqXbZKcuJE+GQT7/0/E9+Rcun4Cu3tiqKIZU62IVpNZhOsSbgJEc44GvsyPt1
tSjJ7Idk+MAFOgOTJQznzHTHi5o3LMADlRZGWEykt/chuwWEATQ9jqvW8ZMbKN5XpjJ3UyIN4GcK
IKRiUxOPBeyjXvwVqM1mYipyKtENqWmlKFTwfUu98iNY7mrvCd3lTYi0Vd6oCjXXavaRWvSIdDYl
6oRLhmY9K2pWHhGL6cHC6l68Nde1sjR3HTvRRaYtyMOE+2gZ/GYylPjgepxPda9NWj6hzOKbJpw+
UXmKxhdI7DHGDgcXMNvO2KpRv0vJOj+++t44a1BKC61p7lQHT3cdGUMQ663u3RzOj77iODAEmV/O
FziTubFnRF40IRWjHE2Y7+8CVw3RDpE5zduC1UJuPZvrryyDLsS/AKMi7CmZkgth9xm0NPWYlsUP
uCDze45ObOCqYLAynFEwyR4YDGJCgi83VbsUXStnMO96Fty8zvhgjGnz+USrWNK30RL85DmBaoRR
AZXDQ1giVeolKT7c7rQmKjU7JPbWjINOti0nTv5rNuJRS+WX5Bt9qRF+1FoJSSfAH7gTlctBheYo
tE661Ah8GOpDQz6QcWEJoDpfiTFkMCdG8l0NQG5aONHnGuT/KZtuaKv9FTWn6rAJsWZ2R0eWJpHg
pA5KUUWuiKSb7k46h32RFKIIkAknnreNMqBtfM3QY61pogb8lGywbtoOiKJJCExxwTfte1QaRIPF
V2JxZTtcGkwXVT4WtDqWa0XG9wdYeG+ubiRRRjVJBrtr0sLxZ74CmM7WYn0kZKg+H3sFdlnXGsOO
ogbW3KrxTPa6lD/5O1NVuBw6bYlydBP/1sLZ21j9i1n1LS0NdNv+xCreFdCNcgctnXvGhpkPgauM
rLQBv1VwPSpP6AHwn+S697bRA3dWEfnXn7uLCCCswKYtvXItzOph8EynSDQ93JVg4fVSavmI+nJH
6aEkLhvzWDSx2HCfkjULBhEkE1l68z6ndkS4USob06BKPUiQlcRxtYv969JU+j4jQZuzsx5Sg894
DA6Iqt7kfRBTpcY612V0yphUAOnuEzIZz2HAeTRyYExncWRJtIr9g79bwCYWHoWKe2gBlY7VCz7M
TgXlPnJKJzsMI01bgK+RBrhZKDKorLTfxJ3bKe+0+RIcIZivSgwbH9eOPDWKg+u8/QqRnyHWJHG3
IKWdUHEOnQ/bl0pEqpf4KO5zXxTRcqRnUX3SpnNrkBLnxp8tFMP2kZVBzSxyXAW/YDm35mcQWBb5
TM7r43R6r1rutavGNQWkjD/iOT6VXyXL3UR+XOZyqOAAfQnXB0fGwk+Vth0NJNF0gMl746sGEtN8
nbTZi/RGN1DWoyOG2w6CWqrf5NzT/D/apO5WydkyD2aBLoYNvV6hHR5rA5h4AMmybv5ehE4ft+lr
EMXqs6CzwKYcep/2RT3j3/oLTwmsdHBXE7aGLR8UWqG5nJ0z9p+CDCN+mFicvdtB2TfHQQqu2sIx
eBmDkK18f+Ko1iCnQx3eL22MzovH+isyd+hhBCx1U3AxRvKDmK/ABhNEAAMcIMNNA+45lmwJKLNg
BiXIajyYFWm7EwKPAf5yJjAEnylUdu/nJ4Mk/IL4C6wYpTj+hwdSop3myvXGhDLW6/tNQXLCI7zw
Qe0Yi7O+Qk47iLdX8Dt0jdOse7DYjLCGjDa1juh4JF46L0Gtz9/hoHRUscEGIBOy0tIogvFANLZp
hY9zfIhQX0/a20Hl9En6jDwJGptippMir7WKtPfdO0ts9IyHxF34IAnG5qYcdNJBL5t203BRjmBT
uayV1dOqaRYoqb248JHRyJ+biQYm6Vn8o0D/Kq2LeqJw5R6tJMoDL88Xz/jOzqKh0q7LN9MhHuZ0
tOzle+KwZnZnaIMe8Ojs3ofejF3XL2mXl6wg+X0RKvriaTv1JVtyQDzW23Hmq7mW1NV1ktNkrkBo
hn57rBdAK9aspgtSzkmHjQLjbJhAcT00imtXbID1iNbgdiQPOu5S+SAXD3J6A1x22BEOzaz3K2VA
IgUYleFGsdrB7PtpV35uQMWEZGWw/pBxsAskMNSdGd07cXG/CX18xvZcDx2K1Dc03tB5rE3N6vT0
M5V6l8Y8RLxdeZjvIBhMatxgWAzwfxLi8LyVJFV8jTVbirmMa3VXzwLmME1mW81F3Pzo+gfcJc2y
GI+4UiFOWnwtui1sVRqrJJZ0tc7Z7ZftbFMOKz7pbE41p/wqrkQD/gdMA1wb/74j8p4AYN7+A1hJ
JRGwbYqw6qjUM/KQwjb/8oErBDIVdTxDb0zxoI/83qKR9SjZJxLjOE51S/Ci/7yztBPtTzqbs+Ny
F5hmrWR64VjwTrzuhnzD9lE8fJDwJMONJIxxezfZ3kZJp2Q8TWCoCLGLHRmyO4TjAkHrTIwdgXS9
h9oRFgbtItKu12+SLmMfMgyOWeagkE2z3KExaJ01di4CAJHk/IA7GaZ9BRpA7hTIbtH12acD8aBD
VahL1PVMRBewWR2afB9ygOv2ell9WoPnWn/C4BrrxVGJuOrQJUjGw3vZDXQA/f9v/lV3DYhwK3g2
wXC23f8C9DuwrCbGGRGTXYM9OYX1kGiHpfaOi/5gTStgxSiuwj64H93zcoLaZY4JCXGChgy/ecX4
jcl2Kn/f8k/A1BlRkXXRGtOCkknkIfAWfS+jB2LUcycqbTOPJZOGOx0781evbO/I89l6YPtgwQjh
uVn6WBq5cIt0wWl6O8m3zEmsjUqIhm7XPN32ysBNqp8pnv4GGdAVrlV6TqzjeCcDREjMDnWu4y0H
xAlxLomJUfCNzD9xkcYKBmKMT9TjHsM1FVNEAwwDPl4UUwshQuFbt4QikWugEMVf6ODi0owbgPSy
jy5jx3AZSD0ymSBJK24DGFomvm6/3cVeYW5iEGJL2v1+urmDm0JeiH2tcqThDSKlS38K/OEpzmcX
mZs7ceVRfSPtO+CnFJiGuLiSPOGqvGxTdYwdfgBZo3LvcqRDOrBroNMbhneexJnAv/iw1ZGTyGte
Cw5Z3Wb9aNsOyRLJxcUyqJ5Yo5/GtP295lcmeoCB66u3jPWZXo3lx8i8gY8d/Za4nHaSRUCUZCFr
I7VKbq0hMi2+NS8FOAytwugCbbhiDX9pKCmS7owsp5/6Dn6wLWlkHeYz2NOlvQXAHM4tthB0fJbW
Gb4CPUVcBDCXqakh8SciCO/jt9BDCpMp1uJnr7/26ftsYelzWhEGh1WVt6ta99A9bOv/9sr3uBF2
o4igu0onNwdSgxhSrY5ps09YSxoy3CVzWJO1UhQYzmLEsHpJRomauE88Wu+Xux57z4KAjrUfBsrH
Wlwk5ZfMvdJz25D8VzdqRXh1sHblzBQRh93N1/9op3Q5TZ+lbHPsRnoNKBXYxAjWx+rb1+XwYOjq
+Q+3U+h7bladCZ7g+xoebO4vkKHFFIPsE0ct7BmZXIqWhYQCxlCsL2zz2NjerPZQ31WFrWCVUuFF
jqZe0YUKObnvCtw/m6SDwy5Kgd1nOlsEn7y8CUpRL72BP7djcOdsOvm1DzjDzeCxF8Ag2Xjt2lLY
0+P0zBxgWk1n5ODnkSy+9NKTKDTFElGivspEOkb66rLEtLrSGStI6PRHhlz2gBV51C5+Ly2IM8Up
Zd+oDblR7DOZ8hnM17ujjpIGYHofA+tbq3LIE9FLGV/D7OqIeOisY3bynae2v+TEs1ksJN1TlEOJ
uU9kg8PcBkmvfna7ThraE3vs6DemHyQ/0j0IHo1uKwpn5q/90N5vQTO+h0EAuFa4IGpZQ2FFCo3a
bXHsOV5Uwk4QtejM4ZvfFHn3fNLXA10sfbC0MD3dqRDpEFcubG/xPDT6Bin0n9R+CkPfk/54/giY
EwpjL0wwUfGmCvoaSisBVk4ehULkfzWearM1DYt5+qprBSuAM+wsome3niw8UUj5fFjZHuvZYena
igmZnadkZ/1LdcNPO4UfuTErJ+4ymqmO+Yt/ncvBdl7yNN+nrRsPn5gqq43qibvvS6c6ZhYMLQFV
gr1Himz1haTwDyQdfRcFGGDDj53wz3YDYierFHenA1LSctWPl3Bnsz2zlnn67YrJHUXIGB6SHtJs
snNJtVqdVF3Pc9Qy1h9X6x+znalc2OjOFbe+XpUCxIqrcmYgFbP+xhC/M85eze5JyNEX4dpq1zNS
uuli2W24UEMvLjPimnrOYYAnU+sjQFgjJFifC9p7Nx/a+GNWOntUy4ar/Ci0YsJDdwZ7dx8hzQjD
f6ubGgdy0j9w4H9iWrLbo8CoerdB8nk6OE1oKQTKIH4RcN50pZyT7yt5WmXadquXaPY25GJM1rnY
i7F+qUmP2gA5DNL6aYaVRX80C6kw15aTZQbbO8C3TS8qns6gMf9Dzlv+dsEgDwcOrWdJs45U8U2K
rCmGQNdR0Z7uolXALTuy9w6YwGHlhHcEVOCPf3IfSE37/6wraeZ81wK97VOz7MTsOfL8FqHSaJRX
u2kmyav7wu7bMduCjWmwo7/7ZcbgjfQQUKOY67eN0965UhegfwSqHZGoRwDOOK5+diwyEUbALtBY
V1Pr9xvlQjKSf/KDc3uid6STQ/BTHPWvqTqlPguCNekbc7932IfcSmX2H5JexBV+ho8AjNQ5Uoqy
h1x1VqGMvDcr+LQ+YL0++/AZ7qzWksdIR/gsnzyuYRb7RnjEiuLP5Ga8uq+zLOuehc+CqjH0uk17
RS3DkoxgmXumyEcVZyRqJO6zPFbD5jX5QNJEI1XTdUyv1GHWwd2MtT8MaYsUnkWkzkf6Q7MV1XzI
HmfM/38neZxLIwnjX2///ZLMxKHL3QO0cjlCH6kwOedasFYkFTI1zcTEq7CQyp3YnSsTiRVcQ74M
FR5TurFL7MKXjcWEkqV566jP2yApjPMI4rDmTz2wf3S8X4U9rWq+mcVEehHPgSkrFMNUp6EjNbxw
OmeQImfdG1XvI/aC3K9VTMGlwI0fnqTRaJNH6Oe5sPWZXVNg7Jb0BlnvrAjztALWq8cTVY2iTl9U
BEVdTjlf689z8CzS9WIKNshLd75Hr5KCXQSMitg/V/HR0nRtRkAed/ekC/uXKe6jfoM5HSg3+VhF
ksO4y6e2fJB4UlbycsgiWDJd4NPpTzR5DcZVpzgIjEMCmbM2B1yp5GFiJJk3YBJj9y4ZUKGSnmiD
LpTGNgRaQP2Ia50G8ic1IZs80dZdnbJs8WkpJ0XKH7jVy1v4WNw8tPhxh1vejVe10MqDySXIOmlW
ghEqgmsiPYhDW5Ny7kdipSly3W3Mk+znN4zQ3wHvfugH+6jsyRxKqGCaXIlCcR6sdZCmiaYzOaEs
aekjxozMLuOlClHIkhYI8TEpyXvOSixD2Rc0pPrkCVEhV65AISdhm1NxYJXVeH/n4+uixuDRpEuF
JeWoY3Dw3l9niQZ4O8OhJMdl4U7te/6WQmznnsilYFPqXM1D+DbW8G6GDPb+7EyT1S4qyE7wY7r8
rpQotGRgLRREho1FYEjysm3b6XAqknvM/wRIjo7S2UzVa9jiLCOKlqhyRyTdmWjL5a6bs9WyLReT
sidllqrYiRGFtADR3WvHlmjiNAuloEWpmLt88w/3WBY8xAnO0Fri/srEvjEwTWrGcqSnlM10WkF0
hzi7GVdLM77md2Ss52nNMgBoaj7zlNL4zwM5PIYWwOYcQDpH27G4Z7GwxQyvRIbeeSkHKJ5ZPmdy
7/WdsToOnxt3FaRhrxVEmaHBsczz92x4LCRwvdTYJRi+1Ke4VUtxJxxVSJZJksSNOKU/bmJ7JthM
EsSBZgG95fJzJurl/20N30o7w9fF9V0GytKhgatdSty1QDVb5t8naH4CnakhRzZWYBd3Hec0YNoV
WrKkyEfjeNAj9haGxn5Lhl1sDAlP2bP3lHJFwnwgmtVb07S4fYJzqDp7BlYPnDPSADB9fdUAswsv
D1OV6kilYR5TOPkGoWYuMDOCrJnIWyko0yTkNnbbwVyViuw2NViKCfsFm1D9A3xK6dHCyhOL5Sxo
VpHfhtLqMW1ruYh3WEsccQv/7ZKjHIdBZ+cejCMvlr2LV+Msw934nUDM26V5TMtJ7QQgeBpLDihm
8v/p0cmRbTzKyRMjNhcHvWeUTLvu7qkTAKSBNJAaiMDqc3fk+OvnZ5NJv+J5B+P2uUC+aiCggeRz
TRBI7dpMDBVJsgroKITwVrG3fDXUJxJUhiVIm3dK9SyY82o2ilDUncnL6MgWpvj3h+G+Ws+gMAFn
zKfO/SMBSKF+gbUKBgwSOgdSCFaXIv81MFt5Pi/wRHykVCoB4a851jlf7ySAlIhEmNhIJOrJ2RC1
+iWAkWcYuj+QYGtanAQczv4QThWs923ryK46IfO5Qrdw++1GS7UB7gpqPs1oUMY3IdgcbD+xFjxz
4wxOge29nXiNLMb4YwjbOm044cVodMI84UgAMbBKwahLuCb3lrfXIWjGt3HuPtuDE0KBiS9DgqNo
/Ue2EGaGaZlhjnPSIYY92lJ5J5lIvIuY4UQeLEmsOvnUosTNU9bZ+kNE1GMiMFwXWwnJ6Rdv3Zdz
CrkeJUaaUsG0TGRay7N2czQffJMFU0dnS3PWPSBfyFEP9qA7bnORjjyOSvrecu52CZoFjWprHrsT
Y1lCezqju+i8g0fgzzSOV+SvEqMnPybjD43fTw2+7DH2XwcPq8VIQ/NLtK9juRGcvbDOVNLYYD73
jr5J6OraghTqzIAJ3pCBKsgMtOUe55XpRJU+tpRICtPYiSlgxCIQvppckF9pzNQrQbbp/9VSRAZw
D2VwWsj9lSj8PvQt5kuU/n11XVRSvd67tc+VDEWOEKxKNt+V8/OMllTilZejhGH90zm/1TSTjA2h
R0q0tDlLNDMwlukK+P2KDQCFs0jN7HtUl7WvJmLY+Zm3O7eMs/NMLnjXylM3xfCyIwgmDyRJZ0uo
YZwdCMSnIWhzld//5jZSxo0DtzjMEJq6Y9VeWlIgHEht5o+yJoK3Kl4SpmdVn1ViXSNkPCE7csnI
2PrkEu9nGhKJsMluXtSpANeB1CGnWhcaMwq4sSDgJP9zShGgu/bK/QQNeoqerLh4xXbXCXgK9zQR
zCX5dMocDYnAwqHS7b34KKA2qMufNjl+bNgexo7vKIh+OvWcD7Rh5NJaGBHhrrbyhTPw3ihFnYvV
3VYC9+QrJlpeBDXScFg2ZcNK7f/gCRt6ykHD1QAbJdBu1PlkMbqJG1IPXbyyJ7/y48bwhj4rysyI
TrOWk3/3hF9I2HB/4qc1yZz/APuo2UiBU81AakQh0Zm2rIdm8L3d+IBGBvyWAmLK1YlvL4NMcH20
Jdd8aIrghyU3edayy9LU5YOIkCdUXMjfaSkrXJFjD7lJkIunkdVwlriAc2fwH2A9PZdn0ck5bMFX
UnWGwPoHPHlbEW+LIPJS5gjbtnQhxlcE5R1ecJBxgwKo2coFwPy6sAsiKG6/72xgMiB9xry70PA+
iViuGrQs+jlfz7AJjy3Sv+8d33OmL0qC7bLwlkGf0edgs4b3rn8aWuqr6dEIOw4J42X6sjd49Z4S
rIXR7dcjY0jjrnRK3TJhniKsnMsz27x368BUY/rThfwl/a/JnoMF6/jyUp5SJyE1Q+kUCx1QNQPJ
3I7Hd6BPsjTwelDCTjpFFm0Y/tXgVscYDJQpU+bUH+ezmYvAYppBmiSFxoED11rD0yxiFZz28jr/
rDTF5Iue8AwR3dGC4BouyTX/MdS+M94mIvOGRt3TLY72EjpOl05QMVFnYDXCPWWAQQrBGTMDXJD8
qSIYhGJeZb+CLQ/PCxlvg4c5wE3Zu4DnZrG5qH0zj79WyFGRw4Fry/Ckz4mGMPmxKIQ6fxs//Fqx
xMcis6Te5RSVhOzl497u3gpV553V+a1FEHcrPIW5nfyAQteYsS1RN/UPGal0iES8WdEUAtpGTqDB
s1UHLYRf96jhjTzcn99zkT5DnyJEScDJup53jDGwDF+zVbAKAz/jKbbqguGe3jhScIGWn5l1/GGe
FvQRJp2O7tOiVO+POLqLWxfFVx0/uKgJEQb6pkwSGS2MG6DXKg/bgUAX/NcDLfjflXpQtj7bBUpV
/hlNcNjb1zVTEHAnXYwssaVZ928/8GLNK2EkPX5FZ7PEOrgbIN/tNkbMqqxnzLDnILwEJoltC7Pt
9bZd/rOuTjBafXBk4ksLmYMgX1oCrCKBuGoN/uRckDyWkL0Xi3j522JJjvl308gLeozKPA+Ttge4
igneYac7Jr+lUfeWoOMyq2zVML1kXeTIhjoswDiGhAC6aDPza3CHMGfpME3crpRxj1dxFQubZXUJ
Ej+EGK40hUryjeT71235FnTHlsghUdSRR7QqmamJYUqxyJfIBP+9FSaREPrRYxvNBQHsmpgM2JEH
f6zx8D1mHQ/QoWn9BuCO47OBGRky/8B7erlEAhCqIQee5t4GB8ZJnlXBAjNq2Vst21DIVwFlay8k
NGuPiP1JHeUvWzWEhepjcj8QNHfqcIc1dCDoTxJcCu3oZP9FNVnIj3l2SH/alDmt4urI4YJkRINo
aLRjXMxCIqqQBCrg8kbCYE24sZbWD5tMn8YGaW+3Rxx0F5C9lnLd80ZQ3H6r9fN9nL+OVIzBuk4P
zHxe4RN7P+levSQT7CGZdcEtYbPzgLRUa0ftxJkn8OUidXxYM1JaXLIWN6BwN/OidY2mKfxuTn9d
Zryau0eu3hrB0VetsDwVbLM5AoWhfuR5a3xzQe3dlJimPb0FqCZwnis5ylujECe8VZ7eH/sU6vn4
B9kTaprMbbGAvNt8sx5272E5H7kArdDwWl1S68unbt5owaswPjVL8z6MNLNHeDM4iBppnBuo17Nh
qjOY/DPowvImQAEuZehsGyN3GfsTRQpeHq/2P+vhHHazHg+QfzBv8N8kv2KFG4J/kd1uJsbsqmew
5IaOwt4XHY2DlNIWXxD8WteIQmfVqfCfu8E5rft4AT08N3sZmQ5vvUr4CN7Xo12WwknX2QcpUCxm
WQggFYQB1HVWOS9nOVCXUFtfZfj/2vFQH3tzjI3NeJ1vUWjKMMbnzLTD+dDwZjFlo6VT/3pBhPxv
wUairb4BWlNXbcVBE7YjQSkymhBD3d8Yc/hdPDENf2uBb/iBkdfUnEphxItZ0K1KLt7YbRqrkCH6
zeWzltcoe4TBjxMoEGsGwSs4NxQpcy+ejCpndYKO5Jq2WJjx9H4bk2Ot2fypim1o16jqSslYD65G
0TMSQcGgugnL90ku1RTcs6aVpGDNHGDhr84DjaDoyRFQs1iP5uuQADvWdijsxEnMOpFUyJ3N5XN+
LTcehZ+otpeNp35sdYKk+tm1KXRc2H8L4Ss82tVsoH86AO/roXU+KiHCC0jE3WF23qAyg9U2fQ37
slHa9DRLd1ig+00bFAaXUXtzhmg7EoP9kCCFGjhotfgICzC7zv4T0BE7yOOfX8K7Sen+KdFTG9Z3
JJBtZJLNiz2LK8mdm7sYfp3af0c5L1c2ZKRMoYfIhFBifq5g7cgKJAmCFbR7bQdP0APMNQjJwLBo
/vE66EuXfo32LfCtwcqQz9PGTvKqXNxX3yFLLqpsEApjnXxNEJoTq57ov3HPESCqrrZ1e6ugDC3p
iKnTCbRfZPW7zJkaNNElGyG6ZpIWtNqm+wuP1gUJsAci4u9U0uNn+eCNiBLQvGhrDSt3Y61Urara
/1m49JlPdLhshHb/Xkn+7QdFuvfFngtUkSX0dAzcbGOaRdlWhOkrwBaAjsOzcJfozVuq4FFWbZil
sGVb8bT+KjxM0hoV6sbjxEpJnCRuKfWUoIIrxqPAXjV0+pUhtVOgCPF1XLVdPdbOgvauFuLne4Fv
9MzlfZpaZj0aN6lTtm4FhCDxU/lrdHgjRBG6LFmXtR6d3un6K2749D6aiHhXhB/xCt0Qu2BTco5G
nrg8lxrc//LPHQw1Bn4FSii9aE0OLlwxw34LvU5xOpFL2Jw85ly1m+4dLBnKk7Zt33X5h0RUjXpa
ji1g91nKKXPNAO9/gr3P47NhjC857Ts8fqwrFlB7k5r20lAN7WV7C3oWAAa5aRtvCEkyw8LtLvH0
8G6lFYNDwwQdcsPnUk3CXU9OLIL6EEnZ5+WJx0gXLdwaSGti3vi7Z8tv+23WHfM8eL1PbyKOeoS+
DNjXb3xgtREgzapwV7fY17r06/fnQOV117ebYymxo7l6HwyxXtmxOZgpjT0FT0nD6JhsA/rkypQM
d5rRmbjrxe97mhTklFsWjCBiP4b2K9Rdsg0/l/HjpP976788AYF1FHyuHKImwBgP0oeWHmAjLQkM
b39q7AamHAjuRT0Rit4Ih5BwIHADAfZ0fKXFPzilMssLquHIjMvAv/U2+5Q0rfga9JHtskeSG26S
SzvDsIcjQ3SHaw+GDMqK8PtvGYuLgxYHeHWZkN3YDGq5k2PEA8Vxm1tBTf7BkD+mWztK1AW3lTna
4N21zp5njz7+TlPQL8EfBZpx207j1T/4yRhGZ34OYDnkE1erjhWz+OPhRxbFvl1hWD2iImcYcpiV
zaJ/Qu6lPO66t32yYMYCJeHiHHSPCzy0vmnALS4UtWlnUDt99Fd3+EEzv4EPnh0376Kzm5LR/Bdj
1/90Shca07DVTYlnYHS2itexOOCjQSmYUELe8oM6YR15JIvvbpn62BRX/EqRyWYDXO6G6XGpLDuf
LHfL6XhPPErjLFm205i7CF232jEUpYytbq9XyMf73EzaS1xXAGpHJg7chNSkFRYBjiMnQIyCUHYx
Y87+JycaiSD6JaBiL2pVVNzJnVqdsHAYqyu4cUi+f91sdC67vNLdxmu8/Bejaokr468pmdez2VaV
vGhgbuXxyZyTi0jL06D4IA8EkB3Q/ZO5BoYAk0DGNplKqeZTOxMQ4M03i+nH49H+hXOy0BQ6N3Sy
1E2CQxDfqD6zVucCDjzKSfz52XJj8GCsFQI14+9wQDKy19rlNmzxq+1F+HxIgaFJtowz2hTIUbHo
96eUUv0NkkKaRJnSmnoBmjCfVAIi0yezUjALOLene/P+iBiq7S35S+Mwv1e2Ube3A0+t3dgweIqV
tM+YGDdlS79Pc0R7dPYm/5iOCUA0Zxj1Iuy2QFRbV3OEpmo2SMHYeF6x1zUrIsOVoSpiHsZWLRoN
nuCVjrVV/q26Gt8oUqawsnJzwLvyW/jK2vJIdris+3PNde0VfLnI2+Q4qjyj9WQ2865KAa52+xD2
irfgQrwMPucrS44nHRIUsWeTwggflxuVPgrZ2cTsnCbtVX4vXC1ub8+zRCI7iiiexU4dV9rB9xJR
vr52dF6mZOXxG2brwtuj6DX3RotrtkAKI6xLctPNdMoH9TUaObzh8r441C1wNwAKNv/zEBiRMzNE
nvRSqYGsyHV8VL55YZzk2pcqCGGx4358KzdFyjPuWq/3iVrBnRbK7SI7W1+1XGci9++9fuwZARvV
yzCSRzqWSNjlhJChpqnhO6cZvrehKLICjJ+IyWe/4GtDSvosCV3B51bg4mPA7UgV3rP4w2yRKn1C
ZGMj4kkjVJLslt+uEP3jNtxfOzYqtJKBGDQ+iYtM0Nr3jzzTvery/1sm8TNVokj+uSPslpx2QSzF
su3GlbQWj5MWJ81dPenQlyuUxdsRi57C6bwycz5QbtC+Jxma+Vj94JYY7zCw9FIUl+RDqw3pgzMT
pD0fRwhP+YwNvWrqjNt2lp94DzjoTa8DWfVmR22Vmtv1tJjfVHU3p0DEecv1AF+WvIOKx3MhiMI/
SddL6ScpbeWxExhASvZLwj3fdzkUjwIab58vDCn/+Q6NTMJWUiIahYAa6ZHDeTdn7m3Tk82cNyTJ
erVAw9JenC/H4TEBdrLgGiePF4M3mcT7MFtrvc1F0vUtis1nY1xN+B/3IFQC4ACauLOrCVMNz7/l
0jM3eTaCVJ5iTkrWS3uW17BkPxZf9QFtKeSUnKKQMmTWDE0njXHtSQIk/vWbR++gl1kW6iOkK8yZ
bMUhwkXBDJG+J/uVhxsW1FJnw7JQfAFGnh6hNlMrTbSbEY7OmydB0uX35KDrPjPpSbSKyBGlhrOK
sSOTZ9zN1qR2VCT7CiZUyiVbwUsKb9QzSnXZZoWyRW08xWJxuMDFciyZiLDvTlm6k+ymUl5SIB9M
f9yJ93jVPktE/bOyybPTrtIYgvk73Wcf+N4/Du8+PWLK0aI9/TEnqX6N1Lb69+fpd18WRSy9061a
qdNbpTSFinJqKS5mY1Vd9cIh2/y2zzTQ1CEqQEcTDQ65KzWmhHU8vwzo46KBG7u9VYgHO81AAsJO
4gXazHw5owah9l/OF0GqS4bVJCkOfhlfkCpSC1z/CHBtk1H9efv55oAfW0I0QsR/IgTkpfySV/Ie
IUibFQOJPGF3CuiCOZ23nsMNehD+hkwMIsaUE6V8GwR172KmMlyG2BpMztnIxuClrM7yC/nY4YRI
suqTosl22Rowik7DVo7hUKxbiBCWSkXKwhWBbvIP+pe9JxI8HbFPw2zGilgNRZXWSwk3VmcdpVtj
3BvVQihdhcLKgnRndTas/hUeNzFhh0Zyy5jx7oI6XasIrwSqxUBBzIyS4WUTKtjRrwBXgOfqg76r
7FIWPyY7vnSq5pK74mKAux606gKaawrGzHSimclQAZy6rb+j/547R0D9Ujf2gPYQ0POeiG4qLim2
pKe7cX9BCoprPT8ETqmnFg4tGBUPlFZ7Nwn80P1ZxUuO3SOD7P8nxquGOraKckncEBf35c1JtM5L
2rw74A0xWEiDcCx+oVKN9Aq/1VuwzAozBDIQYK6KyTjcx4qWsNXeyyu3vlTr15rWkeTMhlCDd5fV
mISm3VQlqbyqq/HerIsg7vEwv+gqy6+/mR9GENe3GezcFvHF8kHO7cw262GHXJExkDMXMYiWxoVq
V1iSN2bWncqJL2e52YFvhuCfb6RjYkxYzFeeNNhPPHJ+RH3ndgO7W+VskRIk+FbsaVc1EfkS06U4
Hp2O661a9ji0j8P2cGcGZUpc6cUFw3ml1bT5XYzVGaDHP4Ox9gXl/iYbZHrMoRovGINfXIr4aRMB
TG9IZd1b03RsidEKAU9R9NAZU3Nc43HbfIVN4tde0NVoM2au0u/LHJSydL5PNWDP+dyE59T6jSEe
1Pq+QG5uBIWOIqHlCO+hYb+exHW95tdWX1GlgN+sMmWr3fogpiOHerI+SMF7MkTLHomD6OzCRAAH
YAmx4XpgpgI8/HPrBGxeNUMLfIOLR+6PNZSF8G/wU9RwcwfhwN4ndpPfN5lXv1AuNqIgMw2Oy0gL
fmkYHhppoMkBnWMB4miWHS+26HPUjvrhHswEJpKXqiIeP4SKWw3yGdUGSurTPosotkbQU4HCBCUu
DfarbAoiSR7ew/EfYELfiWoJeeHEzDexZUsjyL6ZMFD3dwhKq15L2vBIEnqmP1eBjbfFIB0Ak0lX
j+Cunk60onsc7G2wmRCd8kJgcmcMfSSmidODOk4HjupEP6ELad2JR3hiowmrZ8x3g51O03QUupOH
uzd1VdsGZ/+9gpN1+IrP3a0LFpRWzCgpwk1dX+OycKd/NmJyjy6U63qxuRnvWjltsgzhwFtFfgg9
mq0PRhkFh1fIG7F64nLWPr/u9RK14IT3MhFTRryoqH6aLoSs8W21QgsO/79SN73yY4NEjbXvPwag
fPSmN7FBhX0gbVe5wJSpwyL0/QZcHsVYZnnvYK0LPkuExucTGTMKaU53yLLqtwht9aFm+Y/6pEhO
WqIZziPHq8aqk4BNNLRffD7BlylL6NJYAKsf7zBPwIm6iyInRzAcSaSZ/e2XS5vTYjZvZWrtCjQj
T94vAvSCfNnza2vzs6zwSrVViJ4jXaYDlKey7zQVnS5ZBJoH43dWxdmAkRuUFHq5rem9iC61Dbnw
scJ6znXbGT2s0uAZ170/O1GwClZpqey+MVtFlQeo8WXcKGgny4pWLqJkMo5SDX5LEGc4woEec1B1
Q8kLi4vggl/zqnVpkWrirI6Dgj18GYj8k38SHAc6+3PF0XfQ+CyWyeG+KMDKUqgZKOigOw80gpan
fTXC/Z+fbNNjME0D/a8dTd83glvULz9bJ7JlcjHJ4pHuduv+Pmq5LSRxp2+qhb0EO4H6p4fuNM7X
hBvu0QnKFQO1ZSgFejztPkyDI/IhQcXC4SLLk3MoeONNV45eh/y6PGVmW5PSA2I6o3ovuh6M3saL
WdRsUe1qsX2oJr6z+6FXTziuSqTRcqSZjjoWke+MYj7p5LQiMhSqOdZvSogCU1+mFO4CnhEC68HH
wKvmC366kIA1S4INvp64jf7qvPUzToQnS6eLO74FykHaTRPt5VoO+j9k+GeR25Pg16LUbk/GAdvA
0uuOkfORNyZyCkmImPpOaIBwmsB3bJ979w6nkdBwpgoCDS+F/GLk6oMlF6jZ6RqK7gvs8lYXVmVK
FG0pWNJ10IL51Y0IG3G8/H6M09un7CEsugVtZoTUHlssIuLRSPGLFJZE3IzkYt33xL16iW2RYSuJ
70ll7YXzh1yIPkufnwfASLnwqNbF4Y+9dt+7tg9DrQZgncUGq6qvC45fhl15G38qztAS6tsPEBjL
/+TvfZIoT5pJEHeH3g6TS4RYUFSxXTXD/C+gTuzvN/xY8Rbbi2r1jj77gsMJTFo6ifTuPLyEXWTC
i9w530OAbCfjcnuUCRsoH/24Yc1qQZW55wFou+K7nQgUHYSrNKLOuprlW+OtTMinEN4V0ehExDzn
s7KDjUWS9oMXE43HeTmDp64NODz+UKM9wGHBe0vqPgZqLR7choOQZ8wHQR3WDkwah7VHDnviKUXo
vRLXvBDk0HK/+ZWx0OJO665FggJOls/I/HkRIsdob9C/H1aGJ2PyJx4J7gqRQyb3HwzEn+aw4d5o
hsRUa6GSon0UiwZ2uC8T1NwEo+W8ti6qxTyX/QPHZYuQNP8NvfTuA2embuu6FcWni+fGPbAMG76x
jSHUaWtmkaQyn8YDTs8KB8i9r2TzZ0RNWeAx/SlhZtqAmTo4/7WclhvkEQPQ9C9rtp7cc8tqYYtM
f9mmZPOtU8l4KCuFJgxOPunVjtEk2Z9tlwtwQUwbC6HN375bdli+/9LfHUOZT7Ruyk+/I9+qLPBo
yG/6dS4YiJFmo5/JvVsd1sRsB8O9J0fRZZ7EJLn0rox5kdhzd6/jdALMwje2jPYZlbGQRfrGYDJx
QY3FzuDdVVBH2RRuw2tBUPPMRJhZRg8x6+VwzN4yOnvjCfIV2BTKplSokinoLU2SQ/SvARWBSoFT
EfrAVUgnuD0NnPqANdmJlJY+oY8fVRjAxEo+xZHFS/KweSvpBf/muAPUKiSPxPx0cmFI+AzPA/x/
q+7fQX+PCFZm4J6Bo77qk20sE5vUU197Kv7hnaZOf3msrj1gUljPTDQ0F8iFd1y264oFMtWFlX18
W2AWnu3bVtIcz8yRWqjdKT18qDJ0FqyJofXoSPNiEdfUgfC6OdCT326r4BamHX13eye9KcFSVm8E
2WcQ7cFz2UR4SqslIkXJYdQd55yAPbfxLx0UBbsgXtL5nzpJnktijogGhqh9Yl3M2jQkG6mSRHHu
QhYTn/G+shZpLqoJKpAhczNc6CCpsssCVB+BFwBPo4D1X35Zo+zRHpaDNI6/yIAkskXNAQeJRKah
H9omuSbqMvQzN0Q2pueiR2AmEkuxS5HYnoP1mwUCxhDRZIKv2DXT2D8/9NyPlsvQpYVfWn2j+dyn
+oUdAgGVRbz5grimi8pn3Jk2hYTOR8INETXBlszap8Q4ATEm9ylzHYMOSC1AmnIkFyWZEgrZdlH/
QqZPLtyBm9PYB5bxX39hvfUjfJIYmUzdWxJzT89hkEo0emRfWQmhf8qOEAK0pS81GB1nM0SvR+Zr
x6HQmZ+0cR9NkfK/Te9o+RIbKYkAQAz4rIqEE/HqGAtbSvmdhilpUCdje5W28hinzvjCuXJUuvCQ
CscwZkmGH8dU1mlI0XT6LyEVYDNHaTrFemRtlyMaqhCuRexKGVrPiF2yycusv2+uxtWJp+G4Pyb/
K2S+N1amHMd1kN8H4SMxpCT7z/ks0WDzI8r1KPIqIuqUKaxVX46YQFoozY3LzSzaMxVeytsj69/U
KcgklA1jGdLayBOm++lSyzeFYIFQv91feFkQo9Ot8nyRY23DCFIm512FluyVj+lwTFw3k2hvHdqI
4rLOObd7F/OVRurtgdtCeN8lL0dsSVwqxOnkL2wfoX+nYxAiMWuKQ6ZwA0V92ZmIy9iaer7QZxQu
lat+FpHZmablWDW557++6+BcVIHY5zsD5xfrmrjCtqpTfU701xHg8Gt+a5QM+VbMSeTQ67ucVSkQ
tB6OMt6E3nSuf3pHdl6wITGtv7v87uN91cuRvsHaeP2YZIPbSeceS8dLec9tKGAmb421lyduZ9rx
IPjz2v/4zoCsNYsePaTEpg6ni8wT0dkIAwWP4qHU8NZeR0xyjo+PJGY1Df0qfh4p+P0GPRrjONve
JI28R57iIdaKCWYULiNJI6GkR6qlLqOhH9XafsnSgXnP3VvvQJ62M4/FzroGIn0kDUBIgTtuLZ6U
2UEbKaOxy2I63RozEDAQjJKnYNSyqAu/+n0hvNLvisZzo5Rq4gcbHvHnwcVYjGZaaS+JqPR7MEOh
oVwsIJ0od8R96bR8I8cPIydYbV/gCHbpifIvoHAG5qKqdiqTxcfoy8POoXOO0n1hVvJZex06x6PW
j3STTrp0J1bd0C/Tk53Uw4xyk34MoBeivw4Om7pcuKlW2ERHOAlhb7RJGPugtiq1OqjQkIPpeDCh
BiL2CI5FFgGLl3eircgDksMYnZeL0paKB/a+IQ0fwXbEvkaa2OzjvCxkS4xWxqP0S4biBnVTr/1V
oHIHUcBrW7Xo6wuNvHOv4VDpInpZx4xO+/mmi6Cpc1pKGJhScHBpZeRXiqOQoOyxTpb53a47UNIi
e+6SDmmGH8+lPAScwl0/C45wcyHIemvtOnyIWI+At5Af32MsieeJaw9hRIc7GGaXaikH4TX9XoSx
dcoQgVtpEXzScThg5/ojONv1Q37GEtJ2gZbzQgXdGTGefP3CueSTPbtk2UsZXtVacB5sm9clLwnJ
FbNiB7AJLqCXiyTX6A4XGVPoV7a2Nqsa9tGVN8hVUwpnVjNzQftpzKUixzWV8bxxqd8E4qMqyawc
C23kOPaXjXUhXd/v1WH1KrfE5D1bzBs0dFGnmMHHbcY3Mw43HeASjoHC3V4AWBJNMmdTVihFBD0u
HDuM6AZSaxr+KZKjiaaadEQk8iQJOYYCSCuHiP2zhawgjuJJkLpGbGpEWamXJXKymbDVWOu9X2Kg
Jc9R9M+UugfoEbxbsIotLqXWt2fvaVsHktK1uHSq+5YX5T3IMPyTLeBDYoyjrprO2/2Z/D7fdgrY
u/eZXwI7ruzj8h9DudRgIWtcPMJ0rPa/xRTfLgRQ7TcUPSWMN8cGeO3VozWjgzV3o2l34imHG+PO
4fRh+nKK8aLA/23hgFawHUBRh95gTYMmxrcODEoY9IflRKgLxp235PF5SCBkIkQX2TpNnLoSu70E
JC2JENCfHf5D1b/oZS0n1OXuiJieETmdYWDxyvUSoDxSt5Sn+ASWzK61hKfJyvO+Mdg2kr+PRmQE
qrYMG5bJGU8uEG+qvMPGI/kxBlqaNFMb5b+PPaatojKtr4R6RR32eg5xNoNZPC6cytbAcAmBHYtX
zXWmv1LqIk7ZZmd4P957aBLALIL9ZmbhoP7Xn0rs6hSgzNsh+AdllJglUgK6RCniNN7Mi4sKLX9j
oBPoojO6ktEhQ9F+QyVBmZDCDhuTie78lu5KPc7Jni1k2lRpYUSsEnbXWiJ9Cw+dCtfcgYi3+gBX
VzGta8wR0bQ7BuIx0x2vsjqFFO61M0CpMIy1Oj6imgbesTAFzYSwvMZfj+qfW0CJC2g27lE7+Bh/
02AxhByMOcLElUtHrREffOiuMvQujCwfKsUNYORb7KqY017X51W5WJieKJxMfyAPM9YtFtB7dah9
QN3Ac/j13MobegKgYvv1eeIInrh1/hY99PVSF+oepcwMkgC1zTUaydmtwSDbXfF42r9Q693DWbUg
eHv4bVmVJmpf0peOyZIKCAfgjP91XYgkoA0PolWst3WF56TjqIrU7ZJcg9/TZfj3lhaYtg4tFdiZ
yoL0KZNq56KnpIKNFobWEX5Hd6dpauPIwik8CUn/vq1K6zdda0Quo1gs7xCiLr64gGS7k4IALlb4
Slq626hd0bQ7wSqH2XEKp6WAADjHmx7KT49HipUhxxSOzGkx597Vc+mt3c7QoI4pYmETzYw0GUVe
65m3TNwCWr1shdwZ6LxZrfpeznAxUkFTJb6gEc/reTswRFcbmcPa6LDXU1ef8OTbu6ekYydkCpVM
YNP2HiTXfCgSpeFD5Ij/bmWG11OfYdGaKl9WCDZ517qQgtZwKJzDszxRc0vKn+64zyuqvD6ZNpZQ
NScPFmimXjrP+2lFC7S6mEedLV3sssOP+xzOIiqwTFn/grAMLxVtG2cP5VzXf51F6GmWAXmli6oV
bxWBIfdr3Ua/NyNvdUfppTUv4IUKU/k3hMWw5u/rlYz/i5FpzetsWoni/dQcxhed9vffsR1Z2bmA
mmf8C4Z8rdrdOYP9X7up3e7KFraGc860i1OAc1ifBJooTMY/RkssDmMJoLxQo5+MOpY4IqzWsdPF
auR4/GZ/M8heK2TmJqYMx/5l1MB7jyb6gqMHqBB7eCaKNJXu76Vc60oJhKB7Bi4UyVUCkfUkre6C
vUfl7wBHDv0Gv+sJ/rhfc26KOuRBht092V+knRDNSj0sNfIxm99Ehhd7qYhUo/VzUm6vCeicGksV
WlXzXBOrU6lM6DlSZEyQ88KmEvGbP3Ko7Jx+zw7TQL9bHHzJlkusiyin+IM/CNmQFI0ZBtfnnqDQ
TxImcauCFjeMKSlJ1kw5aVQRbILKJlttLvnHBwjPbEEFLiulBTvFjvj+GIfFDghQzTCeZhZyUznk
aJz5gq3wVAgcpGEpCxBTMeJxMSNfGmuOFLnzIgDzluylfr9LyISxjlovQPHVhqLgIOUE8lywhYQK
HI3mtBQIgdEezirbFBjqs9VbY1FiMLxUVNeo3jHUfD3azJO30DMPyrjtnjNA8xSiCSK8q8j1b7ls
RHL5ZNrj/T8A8bU0kZ8P6tZyhN6KLPa1/ZNCWqjixHBqg2FRfgcEwM+r7Cn7Ii2oaYThsvGckRC3
Q1Vuyl0OPzxYdJYJjaLnoM74+mOeBH4lV7WhbvuAPDRMVay1UU9ngyWdL59TQLbUUiKYad01t071
20+pDm6UHXaRvx6aFHQMOsi9F3OC8DBxyFM7mvCBu470bYy+ElC0l8Um8x/kUwSpSBE/uSJqJGah
XNEOKNrvhc6NH8TYLvIRQvyHbGGirVo+FcYilAdAE9CJivs6HRk5MFmNPnJhXlDopnr1sxLkwVYA
TPL+sCjLHxmX+BosajnNPhA2rBJ87kYK0iw1oLpBHhEXoWeixk65jE+QuEzoUElSzFxJ3ldi7vqJ
Ug7yMH4iojKKYaLpdrW/7D4LZ0SZw7ALHR49CTRMVmnfkKjXj3L4FhU1j1U0HbG6QqSVCj3xVS5X
wwiuVpNEf5V+ZB7WYPSyHmyKvnQxN69Q7VUsZcjlovAPq5mpmwCp648ixpy7VOy6lngKPNejFASl
y9HOCZZq77Lg3f9wds6cMgpF29SwJm5hi/5zt3GS6L4hwUjBMVUPxFJrenDis1m3d5GTIe+H369P
PAfmmP/7zJNuo53YiGeQWPB4OgyRjhNQe7BHoS2jughOEVuOuTT0N9zxx/oeOUXpYfSKTS5T8kIB
0IP6LRq/tiXFbvYueWPvQfZ8d1FzzKB7nALfd1Mnp0M4Op2Z2UQcLpbqqoEeaALWcvqDBk+2ABKv
znes9D9bIm29pOI8igWNJpyjkmJFq0sESN9RNv9P+iozJn+cgaJo/4u13jJcsrzK5FMlXrhQZwFD
TdDkjPJLjhVuAe0/RA8rQdlupjHDOpT3YTjb77ruNR1AiZon64tMgJE02yjzetyTZbrrxe2Yz76t
nWqy/DFRTPQtSK9NRnQGrICRpI4Ff4wBVQUNcaWv5Lwtx24Mda2YSHELo5A0kUEFihzxtKeGQBbi
m+ZCMZ6Yl8lF6bEBEXibSw7w1J4OqTBZV18HghpskD2jDWP8j32q6nqlc0wiusGiRIAh3DQwFKyp
v8TBaR+aF+RTYMPo58RxjwCMfxPSily0CAcAie6fV/CYqVIs8lnkCiC0H3sxHYIH8Qhjef/R6bIF
lp+crv8ZpT25APe+HY6f7DrqGyO5DJKGXYHbd2iBVjPEoz7yIl2EXWAMmqq2r1Tz9Evv52d1EZ1+
gfhtANl9eYBXLjqr3FbPfz9S+INSZXMkAgKGF1YTMEXEsG2XVFp6XS3OQKFVUtZPyC5LIHZtyd3L
3ZGEBVNcto6HDDH7y2eyuNeggsTLZTQ1uTclXDelGi+9aPOeqE+nSc8v7w6S+ASeWK1lt8OfbpFA
J17409uuuPoMo2Cp86j4Bw7HgzTlRr8eUzbMVQ5KONQQ8ALrc5zBqFszDNdTEUkF7ke4MNvpWa1v
4E6VUvYUTEu85fNCKL7CxkWRV63LQLY31E68TwkRXkUsNmwu1EV2He0hODxenql5B44B0Owapf3u
74ZPFQF1cXMjiB6MzhE82qzHmBUI/vc9klJlz2j0KE23Gq05ZEA/iDgzn+JuTGEe/P4KQ+XhTSAe
ZVO++UuGwxqmNLtEYLNycAc0FMYDtOOLvMspSQeLRODlw/l+TiPobDEqaoHHtU665okms0vxBPm+
vvpqTGSvj/boX6LzhTo/QUv+ROTM7Txt2yjmz/LyePAakjU6Gh3vO+qnx8OuOFjm83Qn+oZWzMr4
5E3reC7lxlSp+cEghSxTBvB4KtDEiaKm2/KHelkq4sey50n1gzkybgB5N7k8eA4ALHuLxwR5aF7M
ffQpouxLSfQYb7e8M7Fd9cclQOUJfkrVCmP9kzGrpUQy7UgNrQdHu6M4MlNu5YeMG9YWdkmsl6MT
wG0NJGSlwMZq5qImStOMY08nzjSEA0Lxd8xBQ1D2GRJIMjse+EJt64mdggsDU4Ai6N5dRg9sf8Lq
W3YgUYM8F4JVYqiVKUZDiQ55GUvrwBxRnpqbogUSVIVCaDhDZU+YboU1HP6hlwEYGofZJmCMXNEB
rHDSEjAlW2suXx4WJThNGDeqsKqeyAnsBOZiq73EY3OR71r7/ClXOb7o19yFPKg1IoEhCprKmXKL
RHB19DeXkGVgYb2/+90HeRzhoPNURyNL48rTF+SA3tsb5tAfNpjYmWxFWo9+9cHX7KDB9sh9mAGu
Oc6rr84mDYSeBdrCRDMxYZ4PmLSztYXUBsLLQbJX6PxvZcLiulI8QRFUyaEwJSExP4KKVTfL6TsM
5EXyQhsRxMtyO9bdMWtwKDLJWqSVbui8SC7JPo0eexxOra/9/GUqPCvG23Ym5Uz5t854EZRnxfZF
tgpb0LthcA7qyEwq5F62aoC/J+6ZFTQS88haov5GQbvE+q+wYpqU+1qYh4KT+GT0UVRlSdcQWMBJ
JU0r8rKflss8X5ySnPOuGEhyb3vWjBmLdEchxiXpIWY/crN8ozX6pzJqd5teujDahqZJ7pZbeRjM
bhIt7SwkjEiONoJFrQgbv44DRUml3EYsPV6fc5JyLBLyO4xeHim3Eoto2Lveacv1Hknkv7UDiVO6
AaNpLfHUYPWGnPb8XUTpsI7CKp7qWfyvdxzmRGAOFk153Dx7DyZ292+rm0jNWwXuevLTjoy8vwSI
70fnl2GzR3uAMaUTqEvt5ZVBCIzTCnbQKPG+swtFl/Y0+b/rFBloEQzcFvCNobCK06mGyXSrt5VR
UAJjj4okbnSDR0e0ZBM45wwnCY2Eo5J6AeQiR2m6Zever+3Andyrm+r3al7D2NKGjnofUXhbD0v6
x5zNQD/kmfF+Bqu0WxdvjYg0nUW7G8+/Vm6gVt1oyshLuVim5BIVpRhtph4DhhGz/QiaHIrMMukN
vVyV+deFMGdz8RgAHI28aDFyFFIQ7zAInquf3xI6ZyTCkOY6f53rHWo/EEkdH0GNe9nPovm00KvE
mWgZc0iGX1W5K94OmzqQG0emP2TIQHXQk25wAPIKQkn1xMPBS+S8IAZ7+EQGM/HuccidmSmc6CVN
cyefciIoXiHBKYfcJ0DovxKVSyIEELzrX8cgb/vNLz9xUbE5GcpTJaKhnIMFx5Cgq4+qh41pymsl
evo0wcZgeZ8dhQZtdkYa61cEhBUr1tbCdV2cMxsrFRG84WiCqyNN1cW2zKfixPVXEYItFCSSArYZ
z3LFCnyh9SQyNp3MDKtiRWECUuWKsr/xuAXKc0ab9BvmZo19KQU/fQJ1M5FtRoYQUrvKMY53L1l1
uEE00EiUXe9LH/kh7SIfcK5TkjHpSM4BA8+4poDhm+Cjn1VbEhh/nBZKxlNKqHaaa3BrlhE5xTG2
3EBiF/hGLxlO2c6ZMHUu+pmJpu5wGqflPp92uMzwDdviRIpWK3YPwvm4IztNF14Ft4NtX6SxTtsZ
Sg0sNiN4e+Zeg76zg+BP04Om+GgPXe8CBzEUFJISxmHuWjiWparns0bdQLRUpL1RkgYCiNaXfNzm
lQkBQ3+J42RUGkgb6v3hGRGznL6KjCczoJ5JNhczkqnvCNKYRdc2qG/WXlSrijJyz/vMq9t9+b+M
mV6QOcpQ5KXk8p+gs/I4PY5qDWs8B8ozLuAlI7cEEDsJ4waBDGzkbxDTnJCHQgjwte2Q7gKq1NM6
jzgyIvezKHh1KnonMTjpK9BMjWwaNHNJwaas5IyjyDPWR88Fozh9WUcjJL0JmbC5Zcs2cNvVujog
YKqGgkyu2fIMgG5N8VtISnTbP0L2jaGR9svkEC61pyR1K6qtfHvnthMsXCPOh6kLjD0xe6sawQi9
9z3i1kXAq0pmQ+410So7d++oTVIYDN0Mk+huGHQOMQ/1iDhXr1YJvmY2jxbB2TpCFMQN2MchIh5l
c6IqSxEUhYhzKTrD0Ec+tLiQ2xvwF2aOeBjT3guvUp+VSwSjGDzDnKUQX8CI1mlf39qbzvDKyyev
ARrpd8wzlPQVFkksDLEXI9lSLCR8kSMbeRG0h8WcpaLp/Tpy8KYGAKhShTKjKMC9X4ZM/GEM86ri
oLrzx71PsyDWxKANFKrGXbzTcy9qfrrNBbz1bWDhIjBe8KqJxW+dMy96eNREII6EWzFlMOuXisFh
0dmBI+aPgcaQoIx33+X/AcerSM5A/JwtA9T+gIzdJS1An5oWJmGWK1woWxlZOvd5EGoA/x15bfD/
79w7+0+VTQ6BMcrDiRhIKb2W+mSaF6VPlIb5c2Bk56LMbFgz+i9gu9UQN4dhdo2dQUg0oq7iSJAQ
+oIIbmIroQDk9HMJnIvl7q/zvFTLP8tHkgfROYuTx9vJV6/E2F1aRIWRYjdkALa45cyB4q+5COZc
ZGqwbWBj5neK4qwgajqp1TfU3gmlhBxltcR1U7YZru3bHbBnasKPxjY4WDfJ/3gL6AH1X4ynTV0z
uslxh4/T3dav3TLRg9MIeBpy0gtz40k4tKXg5Yt1zVoKDQ6ZkGiIsW1HE0uMLi1CN7rVSVsmfAAU
cSx6NQZX8P4kIt0T1C1BhrO/Ku9CVln1EWSPJKFSXKrqHQUZmLj+7womyFCedBe/v5ZfjXhfB5SK
uIMrWdXaSeSQLwnU/j80LBBqRUywR7JFuTdIqDYk1lqx0v0NoRUy41+0Twnq3kcQwXnd1zBUxHk1
r24kBqUerPGp8i/myECd5NtuD8SRUJmKTuw77vR6Xkm8AOll22ST9t5d9Gs/r1G///lkDqrVWxpe
Nc9/odzijAPK6R9qpgksnAowgASJbTikIBugGCZhbHP+sQiL9K9WheJEJzm2Wesp/LB/EyceTvlb
oa1EthL+96vnvFyuZSTZ4obyujP6h/w+gQIMTI/SFI/ub9plXaS7t9mxnW/Ue0q8ucHIYIUfoSAS
AutuKe/BjcQV5QvFZ/cQyQJMsJ/KgWaKr6vIh7F6fCSrV8sIk116z0p+VySefJ2uXVnOFTrFt9VH
cBGkNAcQZBPIZJlVNHMcygojYW0ms1mPvCwhj8nV9mCDIYEaaceI1c7qVCgp5x4BOhbfkKTyAJtl
8V8VLVG/kDriUIOBBq7epwA9giOPFwWV5JyOHtXC8D/WUtiIxNh2blTl47WMLElPHB85XbuavV0n
CrjtSaEKBh4PCub82P0amUACIpfILN5MXqzesSZCwQqdQVd3gQuX5TfUzS0iBGlKgsDpXVnbVHbH
SSEtmvksBsytnqMEZGc1z2MGPv9E1xN6EddLEyY/B4s/lQcYkmu6jhbVST33L94M44IWWEAZ2WjP
22eYU/YKuT2HitTedVkwDurhZPKUM1A7yZUv1XuRRSV5/uXJnxQmVClcDuR38Sa59Wq3AJBOPwbn
eYMxLZqC9aW+s1hE78HM24GnEr+y+r3+q2xnf0th7dc4DTlORdUzkeHXn1TbflCpnfcgdw12lNio
RcqNyggI/M1rdErV63gf6c1TUKnnOyjIEQxjphRpIFg/F6b5RjVCzDn9XPOSYTiNTU1/atBLEXYW
BrSMYi25e8I7YStBYXTpqzT++4pK6hmu4QXSzILVJ1z5NCMPvxEFiKooOPh99mmIriAUpqcZqP+u
/K5xMAhMYjFwazKwtUrBBA2UVKei8ZibBmLjQh4vK5XakvV81jm24MW1FTQC+FL6WCoQmgKOOkLj
ynCXl6Md93G6N/Tr2wmptVODk3cvqoPXvd8FGNSv+fx8bNshfY06SJGarBRZIiBCwhqvlo0sIww6
/f139oGHBDx4+PZje/nb9WDbj76zuVvqtOQUa1k4b36xUqOzMQ/OCxEWHR6PJWTu3xMZoWdhWdgz
2sLVXInxRVybT79ufGtWlfIHOo7uiQznkj+0wbB9ECMO2XtJvcftuff0KAUXgT0CGNriEb3lSsUz
wG2tLNd8puyOyTg02pBPI23WxKcVKuFr41iekbOOgAcOPSyv8e8apqHllgFzIWMTByxN2GICYom8
oy+kab8WZE+IzjbTt/fDmuZ0o4ZvTQAxluUDjtlvLISY5QAxmlEEcWH6BXerpxHNnIaXLIBX7W5u
JuOTKtWKEgIiigmRmCqdqyGHovCEoiOJ4dP2gZd3SdfXVTQdLUTXA0YGd3a+WB41ID2uNVgelqTe
quRhslqP6oNhpWZjAiuuoJtCsQ/9R6tmmdTN+4TH4eRZwZuKuceBFJIF195JFlD7DMberz5/qKIa
gey54FNn9aRBqG2y3eyyXFCKO2J+pykbRvnPz8kK0TRn3BlSmw8pCEjE8dbLuuoXBSvPClfgPSFO
zGlTedWaIpnrZa4Ru5w1es1GX87LySHEuC8q+ITzoencH2ihKFHxDVJx0eXjCPSouyb69/IgkpEw
w5FHrFQtn9x/FrtCuy6JrocY4j79Kb5V4Xqq9glNXblolzNz76P1I9VOOQO2ijaJKjArYe3h9lYL
Y/oIv4javMeXwHoIBnAGVf9BdnRlWULUpbDvVw8EoJfVkyeuo5jkmyFmOpJErnpw4RVD6VBL+2de
lro18GaKUE7YCniVHpC++mbQI1+aUV0usWO+V97brNAeWITQrPD7NCIHPYITficdwBJyLdmShH/M
8TrhF8AoO+II31oj1gu0R7xPwC0YJh20GvBVx3aCIjHyhfYRiSXHdUyun8MOinFkVnFynPBUeVN8
ZTqudD7zaIieQOa6yxZBYULrorm744R1ZKmcMGda/STxgDHWbeq0DCRfxuYcZSD6g4iJ1M3RQbOf
s8AJ+LYNohFesvR9KVNS4SEDBQxhvZ/D2RVTzgWzlbMfR1ZOoPfwdaRAl6AuWGm9wRjBz1qgGpp9
a/pN7V2CLPZvFw370d3NhM1u57RUjZ0OXu/rpc8+HwfA8+tQekpKShteaQcNIOcZKoHIdjERjFOu
IDVnMV0kwBlMoVHuV5eSmNr2Wmibc+qZd/PRGfnZ4+Ls/D0NfEue7b8bmrVh/yDwL0lBV4sIAKfC
HvwYU9Shgd5XtMibYVYGd042UI0dNBQAYOPYJwt+DfKTVy2qauNy2goAeUPyGhbxnJay0Pcgdw7t
zSdpeAkUXqYpJa5terM8tyxrJN1cHxP3MZU/7rKLlQNZVRFHsrKRuYOcHOHMA+zcQx32XWDPb66Y
Jv8JN/JZJmkru5Ws+TiwBXV4Qr+451ghreZRAN85ggWOz023pNrShNj495US7On11I+z+GUiOwSd
OgPYpcJH/1SSxNx7jD4iPK4jAncuw4l5yPfqPdmbgeG+HeVK8zM58CHAC4ondh6lNHwFtXpm41eM
VEyW0zBYS80264ScaSoymsnGzVtgFUkfDO55O29irsug8/gyII/D1Hjg8suzaTCzEKotB+Y2SPVG
J/KUUOHgVINZ4K9lzfe4WDoqQd/1S7j6wzGRhsky3AjkKSSL+m9szrZrYWo8PS69PuWLQzNVFn+Y
dhh5VFPAydAV12Ffb18nDiICHQBcuW+cq8Y+g0fyq5WgcocU/LJW32a8hVB2z8OdbYTyMR/90l0n
IWwvWV7+e4p4WgXOCprUMsAVEhe81E2VerAowDfyqzzjXCTUlzgWfdSu1L2tE0MvhnU+nS1YD8sy
9ITLDfHI3oP0Y8r8sccwSe4wpFBPwbDsiOA5sPdyP0FtuM2S+/U9+NYUnzBgbqHVqfZouSb5//DN
j4gPRkHt4VOXC7jGAEo5HzBu6m4mClvsNBU00kAzZuVGAOC1VADQ86oW5qNBIM2Dw6M9U6paAXTl
LRxJkToBhLQLT0uwpuZ3QmSb0xUbaq9lm7LcAHDxl+iB7OfekjKJOTiW5AxpgQuajbTpDqjtOTfD
4qZQPd4xPwG4ZIMEo471zYBDPKIBMt8NRyevCXp9pU30SnFfoFxAlumXVhKoXr/jRoNGus4jUB9J
gOT+RreJBA9HuzvDzR+ue2gsLTHNmymx7ucUo7RvWHl58T40jRkUukqSPz4GcCiFPZ3iRp6/lA0q
ZQvKCr8+Nxk/kQ8nbA6ao8vrgov1MmzRCA2QAKXmJhW5piYDumDdVK4Gsb9eCUVI2PDA/6Jl803d
cQCM7xsPUbeHy9ogbL3XglBhoG0/ugJgtBor5qBLyUjLqAhRWxqU7BhWaGDMehm1eLnLMXp7iBBq
+rDo/oTwYSUFsvw0VGvEMIT/G/P7dMUjLr3Q6qdbEvO//MrkomJEDVnV25cJMPqImbYzJ3S4VCPJ
mwXXACh/wHNRAqSleYZrRlazFsMfdI7RSYJUfyC0BRFRfLw+H7hCn7CNS7bq89Yo5UbwAuy+da3T
uaSbzMablF+BIGr2OFLN+z4ymcI3ET3M3H5mjCAzWwioT+vkcRd+GfPxEKtHQD/ZTNVYkjJAzhgk
jAjvfTRerLK0PWNXgjq+0hTw3h8TH+7/U1A6H51hMbwJ2FlFV0cW3u7gGLFb2k16iXQTIw0xkXhs
5l8aSe7WIB7HMFc8EhP08QS1XxeJlTmmFyLQwYxf9NkVF2HWVdVVSuCVIuIMXVBdwsgWkBMoqd0C
E07Y54HRj4kd9yhirC0MULR9RFuxWYaFWCHT1xqVIYJpWHNZQS2MvgONSK1KPKGIbx/DKEd8xwwY
wjatum2ukoY8pG4kwm03TNRqvGetbMWf70UbRSMkT4yhnzRutS+6xpK/mDZ47KFJSi9Vt+F8qp2K
px64OWejhcA0SRJu38xkPMmXEqoxyOv/euHrsta5mdVgRF4UN+G1+FNvUj1KxpIxlznVPevLYGfr
MM4TL8NHLcAceele2caGLJ5I9K/Udm5DX2yT/FZioOqPUuA2ObXZWB0SOylfXAXpSPy18JxQVRay
OVAK1FeZ50WoK27If1Eg1k8FiEhSyb83xOkJiHfHLLsoox7y6zF+ihz8+3N4iiVaesmNni9SwS/D
auqMTncgIdJjPXvjxsxwVQauqzwgF0l3zD2JtXxBx61ZhN7xTOKE2fhkzPGzxwe9gpI9194ylMFJ
3RYNY+Z3lb/3v9tjAfzgAKtsEucjCWD0Az3FIAnWttgTVk41t2vuHFrkQG+j4HUi1+K2Hup3xdeO
UM+hq/VS5gfHf+T0fqv8YappR7el4dtjNgIjMWeTWWLP3+dgY+UtXEixzHidXPAMBbjkiFp+lfuO
fZlT8YrK1lIdjIEf6n9Y5Zo2yHLlIz2Aq5vaVebvN/m2rDWHtnXY+u3DOqNxsG+8dZi/tKwEYq39
A/5+9gpFQ4F8HC7/Z2kAbDNn8gTVedgGNvHXnChDEDPaKBTQHygZND7X2Q/pRMq8vX27jjShJ61E
YjZ4Sh25D/h82avVlcq8JSiMvVjHZWSZeX9MvCA9TCORcCDSZ1AXxa9xMjaMEQ6QGv4UrYkJCs8N
JRlCOPuYvbGwq6xz+egr1pzpUM6NeVHjImmsvYQUnoPX+k6TAyU3DJ2W5LC/wWIVUkZr1lLN15LA
/FUa1t3gkjECzPGySmKg200LLkRR4hvvtETOtJdALxpEFkNQnT6K4+JjIPkt7gy7IgUyir2f+0oo
UShKlWWHYP+cAuMxbBb2UNOS7PFeFEBD8DBxlpoBlu030rmAHoxkxHEah6HbP6y5tyFL9EUbDFy3
kzQHxgLtRcOg71bUQpNNi5fZ6gBoerzBKeECkOmIYo/a48iHwGytPOXJjWuz2PaGnZWCC3/MLXSQ
Nos+lUOpRvYd38DNkDHhjW3GZ0A2HgTzXeC4QeYEpFlSMwmTffeX7UBXR7PBfzItHnUZnwoiosxv
lPlcA/PqQW4RcL/WtIkBM3Seh21hE3E2QswxSHEURvaJeYnkrP7WVq5hYkdxZ+BK0jmXHgF8+GYp
WbQ48pPvnTBTDUzNVyUGlW9RtroFx1KcmF5KzeQi5j/R3wCYMfReIT7NldpFExZrFpU6rhgLhXjd
J3PHcW8Xkxs+dXv41bcG7OCsD0nY7ON1UF/ijPdFNc1YSivGSFmUgljP1IRyD5JLNKgE/nDMOezv
4tQ/Jiqcx8q0Nv5JGQcJPz4xt6A5/Dzx0qJUbudyFN9zuuHO/SjP8xcjx/3jlkSqJ9yONw9eABC/
U1vRlepimHofogbvsVoBnsMslU3JEpp17lgMAh48MpquCjflEU4VJHALR0b1Rc2Ssnj8rF61prt+
OkBR7mBD0+c0xKD9b0mBMSCrT/Gs72kXLgD98/94/VHfF5L8xJVVKu3AUN0yt/gYYDw4ahHWPsFo
QrnL7gBTFIoaaJ1dg1ndKVxNzQtKAGNGHo8CFGEJ4hIFjh00DoCP78v3TNkaVcrp9lU+JrcYUbiQ
GlNzFk1AQFIg20Ol/QAgUEi4BhcDYSuZZVZPqyxNy9dBCH3GpAFVyK7FEeGuLX9W+Kw9hn5Q9Ynp
CciFxI63X4Pgh0RGd0Zr72B73mu5NVJWKeEUbZnJmN1/js+XzK21JfXI/DfV0kSqQnEwQb/Vh6dZ
PYSVlZa9Ur9Me1ymB0J69HKrF91oRQSwogoHEK7honRboF0z9OD5t5qymTnvTmHAkSCTNZRTZO2U
mzUo8fONNz7EfKlOnl6vcs8w0gj+R8TtRAKMlFGVxzbwA8HHZFZXZiocpbtpWVWBZyOWG1yZ/A/6
1D0dGh00PwkRpqSS+tnlf/MNoynTrWCk3Kgnn7V2ub8dVRSRr7y9sp5Ul4mfhSjj2k2CJK2II7Ds
N6WG8hVSg1bwCJF9+vO2VXSYV9N2BWUaE4N/5SbuNydno41KNMH5iZA+Js8AQBsCKoyg+waHQk8O
vTZvRm3n8BW8njopcMopkkozeJfONM+FSvl5NLrb+2WYx521q34gkte8S8HtrHA9TxubFaZzhxIV
YVoNOEnCy2CNMPROstP/d3dpX4DTgfikuQi5zE+FhkNhWroXBWY/umGvxWeqIuhZROmOOMts3wdg
vGxwOuGLPY/sB4NhgUPHSqZ7/ytbA83lDRIHONKrwvkqefzlKkXMzNN0oZmGt8sz3SE3y3rSKaE7
EA/qRNAhXjEgyR2quIBnEoHHF6t6qbZ3KQI7SnZNlu+IvzAPl16JP8Ul/+a5TY/lDopUPIBmGbDi
jbYp+isJhX4e9051R0fAbPgUnZWAuIxsbFNlk3stD1B4LfgA/d49/x5SVwQf+jTMDWohVFVqlRNV
kCqT5qUj7qa0DGLMnvEvdVjNikPXxspXgCNrWMSS/1TebNlCdPT0yTK2Ajk7IjxxRVXy6EVn/G1u
h69uWUjOln0wXtmc3KoDfA4hlbF3Io2svtE6Rvr8zvooqeMXpHZjUOHrZZm6ZvM0QaqSnTLMExJk
OIbzLIFYbSRKE8tmYFTPDFCSLl94RGNJT3ojhx+t10PjkmBxdN+FNMmzB3QI9q2PztBLIOVnauJr
naCtNg0Inu3J26hz2sgfm06f0yRFaRuJQNmN/sTCZgv96W07sPtOmSEoLt0+rz8OdpAmTsdus2OC
juG0rXXZzkT5YzUOjWFERXLtCK2vmejseZKMWnOSS1LqMbMCOfiJ9KWBqrNKFJDXdDLULwRa4nCH
sIHe5rEiFueUWzVdISp0w+17MpmqCtmeWrm6e+EgfPZy/vG7yqm0e9wvKTfTAUWIjpw/V735ktTV
dOnCKVzMfvNS2+ivIEATlq5fFJzHJnWlvc2CzqsRVnyrNWJx/q36VbmEw3xPwRf7/c008niglnAr
lOI5AdjM0tusLX6mqMCisuKRFsy0olt4dtfWMLOoJeNR2DDTQ7VJwG1yRqV7qSlhtXnYqy26RATB
JR5/FI4vd6BiiCrC/0u0IZaQ38MOFxVUZljCS7sQz0z1vWtAlqono3kelKRQAZ9dhcEOXZlZdMbP
qUdBMD/g6CkvERS2HGSLJbNoboWYnV6oLxZ/ZspsvnLsmhSxWPVmv8tka7u6YE4NQmEVHP3ulYWf
Z5wO0HJ12fpJ/+JPRUM/1zzlRL+MpEZI5cAZOsBV1NJYH9gmpFsk58hRnPi7h5MXRqjCMLlBaz8p
SdAhNcfZvBfJn1+6TOqV8+HK0+hn+swDJUgWFlH8cqMUWbnZk0Z/7LAG2O4fxSurzX5dTeqDsF4q
FMIGuK2seMf27wHi9j+OVr7I8wU8f4JzQdW0DAcrbSzeCLROpiDX/FlsHBTSN1Hv+On3hXMNP0+D
ED2sRr0LBN3c9TjaywfeOvNzRhWXJKw0sxH8/yH+VlBKSJWSMEZuBfPuudeDw2DojXyZzA/74eKq
xPRL/mvJqvH3ziIDMi8Vt7mgwBHAmOQ/yVhkcJVm5nI414hRb+HnDjymQj+w7ZeJn3zYWOYvMyxa
3V+sle0s4Ojhk+KZKgC40g9pc0CeiEHqJlvfeYKtsIfwuJpIbCv6CiJb0rgCGW+8pI4J0HYEY1gw
G9vaoxCwZlDtWl87/WA/ZboObhsUtkhjuM4+PgaAf5Qxf4kol10qUdItbhBB8Sz2UMn0xsMlbwAY
LNpl2EJGJXUV4GihK6A9WN4kYQdv3/Etkd+4tJkbbvD6beUcd8YxCylUIoGU6oTR/cl/xEoJ1Q6T
WcSv3HU/EB3g5qEbw0ZRryG4s1Z/A9JarAXLPYAVlTFOajrdg6ir3V3/CYsQ9P6y5oggUSq6z55i
O2O3CRPK0jtmUCqfC3JMQaE9DsTz6aYLd4Clx8FP54mgAOMIY7P9U9ax9P0K4wC4p68KqCdiv8Za
e6wf7qpzWykwCtWNsLhmdSAc6ozZpt0KZErb9pF5t5+pss2ertHrwBDMMVWA4jZTd0F9AkXS1r1p
H4j0F/E+iNLVXGfW6a9l1C9lwyllobsampRP9qzHlfBgkmAK9SUkTekSj3naa2u44cW+wcxCKq70
Kt+ro+H6gkbGJPHGTUJdu5MTgdaJ/B2U9Pr9hxF/9vvaL9gMC47iHu8kcreywa83B16H2/fadACq
3LVWgTIpHzkgPxCTCrW1DLzu7l/wNfA+IQA0euu20+/1+z50TqSm8GY4KYSaTF5KjhslJT/zvnm1
KOsRcssZ/cZUKlABg71eH5wQlqesyT3Ryffhaa/akXfrE/CKU2+9cV4YHpTgUpQtwTvQ040UTow5
EJivdwhPEX+UvaS3vDWjSExV13/dxdZmEGa9PFkas+dwwC9l3Xp8Yrr9uGomHWaFfZ4XCMpmJLtv
48XsugaiDXXIdj2dN1o+A0TgoEFAU2gzacuUVnv56YVKNAGCQMw0Fl+BLtCPcc9oBVDmaZmKRZW3
1tBDHPE7WBh9yJp3Ds+unnl+D7di5eRGRqg7yrzzRKbvIHatnvmheBhLWFExlyuOI+/D0m08d/hd
/u7v2f14bFJV+VOVRqCfIxZkbQvI7pQ6qjP1ypmJ2i/2/Rrw3AfEU4S8MmF2AkCV6v5zUxPhDZnf
H1luH/phpbcdSpneEYA4cBKkdRuGvESvi2cICS2PX/vIpaieulsXqtkKa8kgD3+C9Um0HGfg1jLG
+bElFeKfgN1dsJIRAlpLNQ8njQSh7DFjWmbE9jN+owaM661hAIlBMHjhdkeA7qEchyofjZWCtQEQ
Maoo5pZTPVcqwMbxxfQqwELp8rHKu938+Tv93tbFdrQ/otw6pC1W3LbT6JIWxBgeDgSz3Go6GEhZ
TZznlwWCsNMTF+KSF20Kk3ob0KncNpH0nsDph+w9mpCdNVuLMMyIzafRXLx7V+KfiDmziLHdRaH4
33S04dWrZ7zdtqjvd7CiXZiK2mXGZ4bjBw069xpvjavVQeFvPwydArNV2Il/brwbXu+iZC0wwQle
H9aKl2XQHEPBjlCVKe8Flk2l9GXn9X7LwFmx7Nm8+xNWS9HYRwwMG6ViwJVUeoukAnYejFwcu/AJ
wV7Y0s99tMtxE8TgD1jFLSGDoWGmQbApZFJfAVOj8cVORI5jZMAGEnUYMlMGUCGs6+2B1t5GEXU+
B223YVob5rBBuID76xfPCcHu8FPXKufcYSYQC5eoG7KsgykWKbhD0KxECw5KHh1CMaFgg8Lqrb0d
0i96tMCAMEtw9hCWODgcYc3a2RF6/t+40W+i4zlknQhJGKAPf/ugMnDnHe5Cjyhejsy9Gpj8sRAw
4QnS5LpGsfVvTpAIGCVlSKiK7G7TM+Z6Yq7aYtR14eLk7mz9S31K8miqOIir+UwhlvZ08shoGeBi
DAttqcPiEFkFF+4NlQPmJ74Ovg/lvcTNB+0AKFwS74fWP+DrIw34L1slHZ7D5Wc3XftxgjdLDwPZ
tybzCymDM8a1GvEcV7gJ5If3Lb53LkYgrAUHP97KRtd98ww9cOkawUHh9cM1RYHRPZyJRRSBMp26
0A0ZC6YvZGTc582AEZsdAM0hmY2wrOvt2FzSn26DqpWdlekaXUclbeOtNJA3/O9RWdLH1z1gYi9c
ROjSNBGg8yfOZrFTRdwYVFPFwNWFEB2cUM3QAEyQ5INC8zo5VJPSpz75X6+mNQpo/hl2qLh5nTZb
GzlIAbCEhIJ7XtN0+jiyVwlluug50qzRNaATRqD1uhH6bRL/X+MTzRsF13RtYhZN7mhJxcCgfsVt
JW+3EQMtFzR8nyDHJJkJNGwAAnSGLjstPRfJgR8S7HMnEUtYN7BNORFkX0SMLkAisv1hFaXOUX0c
4aVQJyN700jKkTtE1CHnW6uDa2fn89BFZ4r3IW9K1U+WNZ8iD+BQHsLEl/EdMwB0nvz0c4ca8QwG
cv3j8PkCvLJN5PZ5cHAOXBiE2xgB6/hraMJrkS4k2Wh8og/xYUjCDbHkOyrYnypyJKcX4k0Yc78F
lzR6fbzmgCT89P4foionHnUxnt4F3uN2VYOEfL23+4q1WUUMQ/2K4KA7/KLEb/nw8d6f5E+DXnGV
vR7TLHm6147oM6RlN1tON6chQtsyJ7Rf52DAeEsxIIDc0/2WVtKlmGBFxM5ruwqisAUYmPzNFLvt
O+qCZ2OwUhaQ4OivOqNfeWUF1j4ZZ8q76VG3PqfYdfWB0gTtqGZHYLiAtkQjQuP0UuiMjZJDxEHL
kl3SxeaTmt66b9PaqHREdmhpRxcBcWZLffKhY/9JT/x2oEtZ0Fg594rwWyp0V6Me5EHnJdsuaV26
eyy3SdmkNPi+5ChYBSbsmgRjLEkp6Zobr5Ct4DiEnhD3di+kecfF3A6ZyJ2Ec11ddZz2ZvvXPw4o
megWSDB7Bygw0GVfU9g9mHBltztrBmfXKnSc9midvLsG9eEqP6Z1BY8t7c6r17yLH5e/h2uZKp+2
CkAm6nbTMzYM71UB/KROdlufiCwPmi9j+67CrC3+PkeStwKt8+1mYeqMQTDsnRUUWtO9MnbyVNFk
Ln+fjVH0w2LB3PbEaacL3T3Ls2OCD5Jn4M9T5b8WYGb+/wPKSwpnI98YD0MhKYdXBeJSF8u1U7AC
Ye25uYMoKaTPmsKskfwkkpyP6wz6m380bYGz4AMFLsx6clYDsY7uUJXuJ0h2UcvgYsKDGVuXKh3q
Yy32MTR8atkQ1ao4Wwb9WU90cbe4OGTjf8fmyKd/2dqWgm9EOEelRNHRy9eIzzjkYlx8Gp0ciwd4
ZRhMKqxLhEp/zn7pYZzwYU25z8OMXowD8SWXn1ImbEix+BDOXDH/K7h3jS9mqk811pKy/ly850e4
Tu3uH69G1w7p3KpD8Lx+E5crfzwztamTEI37pCC5JZJ4oETXXyOFj47oxDvrELC7kBCFVV7Z/NS2
EOpcu7BKobh2b7q8bqDnXVaHUai7x3bvQS6nKFQ+UTS1mm+cYOSvbzs+S5CA0boDIWMt5x53z5RC
69XqQurk67KhFLhqxnUIZX19EXTR1/G758h9EFxVx9sT8Mm6/Za1DkSAHFQloQoaRc6hv2YoDSlf
0z+CIWejJCAkb9V0B88DDRQlptIzAJ5s0CF6lnq1nSc1CGMHJ6auEG4Pe6TV9JnB6xSRri/GOjqe
Arah8xEJg9dyXvr/aYJnhKolQYP5Q3lYo+Yjt0TXrT7JGIH8Renf3JnQ4lqvg7ZfCOQg/6WbBDpR
LL+vq24ezTnqLucF3Rf/PCBc6NaxFeYb8bQzCYFlXJHhORw+K1Qe+74PiZIlMcBfEFrGdBvW+eLY
eYRbGiSSGXi5rW7a9MXQbKkZ4UCQWCl6Hfp/fRkRv0Rc40ctfCOsRGDT8eSredH7GmJ22U3I1gU5
FhmcB0H7Mj5MTUYzqA+XIsbcM2gtd7DIiyd7LCmdeVqcT3UmWacp7iK/hKO0gbOEAP5PnQorEND6
vI4ZxaC2hlxNRXE69/uua6e0hubmHs5x+qlxfTL5Xh+OCjPLBznrSpYtuGg1AMt0m/cT0HDuFA1P
8Er3wgfg3DyjSsQm6kAlZy1TWan3/SBOxbGHosa3SLdKrZr/5H3CuveUjFSVZt7trcRm8ol+cC6+
FLDyj6WfcmNgyMf2O2OLR2ZCWSDwaAVZbnYeX/ndypNaXYB2xjImnbmrJ2u6CHhPS1hjytagpHd5
xmWlnuRR8Nh8pNJzSJ7/2m56gC4ohwJpsOyJ2khvkf3uH1d5g1j2f52jttE7VAa8PMFxvjF2Dh3P
xGM9UtSsGbL5yLsLG990TXA2LsiMuLbnefJIzPbzn2dpSmEM4TH+43vecOsVDomaqpxyWV5CnPMS
2lyXeAIthAZMcfhTtp4H2ApkfIxXzA7XdGitgFqhbTGFCNrSEFxrXcw5NWwhnFuJP9IuKyfa7koX
p0ikzoXvXuEcdLmmpvIgfRv+4LoW1sAWn5ZWtv7SyM2VkVjGydguw9ew3b/+np6TpNSpYWeUKnQC
RPrHfym0ZA5ch1GVvqUwaX6djijJn6RD3yMgLpXvcFAY2n7mn84kZNWL3HepI2uTEE0PD1P25c9g
W+1/WAWmJhVZKS9nFJWbq24f6IHBHBOe2J4t4CRZYG9UX1vut4mKJ87FhlVZEU1WrXcPF3WZPnX/
wwsP52u6+8X47hKh5WoHPF+3ptmelnG1reaMBUq9xIzlxOfWdN78tCKR9bBrJnXTkOaCjV8IMx4w
NujTt3zFMg2+ke/j76M3PJ7U+ci4RMZE1uj0KxwHQ4/NhySbc+G5fbl3WH5E5RzEX0v6NDkmXQvr
B7ue2u2J1Kny0RIbg6fRWEek6Vm29YNE33pd3osm20GbXtbxKaLc187aIl7Qs/umLR4iMJqjVxqL
H4UzeATs14G+2SBFbH0LF55F3RYkry55U0zfAHwXB3EaJERNwftmxs98t1lzKyJ62xGHvAgT6tUN
TXQx8YVH+bEbeg8BipU5oXUfMb+hZUL4KfJw0tSg0Z2kih/xM6FOZYxcEiiB4y8pGI5E1hibS4gY
Y6KJoVG0+VXdPAl1rtCJ0XR+S3goPa/uvWqOuuDV5NTrFwfWsLfYder8vjYzrLnTXDC7Qo9xNMgz
BLWgGeuv1NvqjWnisHy4KzFPho5pXJjC75CJUAZ9UeFPYPIfxmZOrziMa8C+lmnnc+QZvvEukGNT
Si1ljFjm6JvCYStR/QTK0ax3v8DoPQiqrZ0+vOmixTXuuRFUrv8ZCilvTPakXtt1Dq8ccgkKLpHM
ZZ61dcnDjm5N9suiVNE5aFpZurJg2laJP81+ZlV2xcAPNC14m3THNybEapLoxYj/So9jAHEHPGrA
KnZeufImHzhvQZQvf28YOMLBLiTuC4g18vnuLF30OhHauMC9jhMzSUwLcNpbk+5f4ajqoNrfbtIU
y5h5E+wpqz86NsznGqNVOATAoW6Vfoie/Hliqv1uQCy4g5hOeIoql/uqRqlN9sPDvy7CltVEHFDN
vCHrxpSwwmuMWD4ELxHX3f0v/5McZ3op4hlcsfwR8LxHG0kXTQvlCkXyRbIY5o1M8OxHDE5OV4cE
WfFh0MdRhG8GUw9bDA9XuA8+Y7c76mdTion4ZE88NzlubrW9EHskQQ1b4Fjon7zjKskWhlFz7Fbl
avIW5Wf69uaPadxVQAMRgltsj7x48lt59YqGYW24YS9imRPX6bLr/+d9CGFtmp4ur4bLs6fXrRUJ
T+1ytYeqdDiUfGxLyNWmODZbY524DgvRgDCXJPtwA2PMtIbDAJpsc+tcFSE4wjHXzpOIqqKbTDtH
A8Ap1fS3mPch+22qo4ZxGvDMXd14EFzMjuAXCvtEouD2IixtnwBnHccNdgEgfqhLXC5qESvWY/4h
JBax0pajXVJ92rzYQBqw0pmS/FP7Hbzxb7Z8/4qPSnuCUtgBskEwrA7LWkVFKGSK5sIUS2Tl7338
hsB7sBFtjJdhN4NY0mBTGt1VPn2X+GHcsuYuIxs/IobT7nMSkQHrCbzWtpItATekoOeJXWVDXq6G
ugmJTUDEjQBS+3Mcn4uH9IX2I/k+tsHq2fCRkrDDTyus6TpHomzHx8EIye2/2PGeQfsuOUF4X2Fh
AsZ5MKtENC8vsp0SjZh9S6Ao1ErpVJ6Wv8AGJXvwbbrGSBVfVaqpov1vkwXLrg5Tze3WkzhJmYZa
f96HHml5Edi0KfZaNpSIURRxjB0fkoEVUv0/NDyEYitpJoTraXjuQ00bNDBLSXAcpj6/mueL/S0h
A3xxdjA5wSNZQf1dCjVfjemH8iLMG9bI/374YAAxTR/M1VV+YxRP822d69NRieNUbED5PaztgrC7
n7kkSbReUhtr6NLoUHYx8s0XkYryKezOIcr15aDw1TZMiwIiaO+VyGJ/5MZg6n+hl37OTDlFc3la
B8EFQhYieJ+GeuGUYaRXFTu7eq+R2nZipy1xY7xtA/kA5+cvhsVPFhS1OlhI00jSzmBaI8w5G2y5
MUia/S1WYBD7RVxHC9SP6puGbPpAzRaFhrZ7cE0Bl2rbzxmf5dDacppTBwpk7S7zpu5PeSnXq7zt
JFj9dEgX3tk4X+DOf2CUTGxEeUC+woyPf5wDoUCwgQlQd121cc8fC88R2E++Nzp5MEUZK5gl7HXn
QItyOWt133rB6ZNQ711Nvb57vZ70IJq1B2dopXWZAEKgYMsOhuYZNnXRMskElY+OpMUT3kYjxHVX
DGNX4pPvuiEuZlKNAFo/DYGT8weNfC7B0Aq7JmEz7yMl6LJn9a/MHv8+9uvmpcH+xR3Hqg/IgdR8
nE36/7MAdJLV+p2LsLNW0Kg7Ig1SYJSeE0ln/Qm7ifaTR8ogBM6GE4IpC+W+cKQU5ycCJnLlhYVp
DJo/R0ar6d+mjNLGlAVJvZ4Vq0Wh4qXq8TELRLdxb4/crL6QeL5E2jjJt3LwUqOyiHxmO/h7h1c0
RUTOItHpFIB/KmDZjF28kIQw6XfVmpwOYC4m3XEhaHaHeiZIYsx+4p40u9zz6qc/I/HqoB3LrgFf
lb6fKF7rHeWbAL/4L3XhdB5OO9tgOBPxf1Y/RRI9kpkbbv3eNlA4IiD1WR5/5r4ro2+gdZCMugC6
2U3oAdbN6zU80OIXmrKmKTOU/5jCg2wOdJ7uTvKTbdBLNQwtJ4zqrHZ8qO6mpPA34j5wFkrGMIZg
80CfjXHtQG2DVwRiC7Y6TDg6xHzcghaR0d8Tv/K7+QLIs/M9LuAwGws/o2R4SVtZ1Nqakzh5L1mU
WKBK/CVDvlt/MyANXy2XPXnYaa63cbxeLS5OVYKbkzKA/p5HfuMA750JCv8skmEmBvFrY9FzDTAa
RkRRad7P3Js8SK5wtKwNTK99mcBz/RaXExWkUTI/T17qLTF7kxwoil4BWsCSg+uMYvjSD5cPDHfz
b3Vrb//zeGze80uaU9oYgM36+s4nlm2phG6Q/Y0eamE0vG3VlRDivAruAeM3oIJQqPjoO0XHAplp
2m16M3NCJoB4EN+m00/Fu/R/wRJBI+r1jv9IAqCGXLaVC7N/INtx5GtvgD3qOVxleqT6E4WRxY3x
yqmYUw21OK+wuSyxKuwzXu+kiEgz2pSvyCCAUL0+TL0AvAdWUWvogJOQHxx5IksAQg2y0G1A/AHZ
tSqpFLM9vfIt9oCBpMPBEKSQc9RcdIUsLe+pgWY0OGBAqzqCg5CxJHB1E8I1U3uOnBbop+GSN/Zz
e5TOqkkouxC8sitd/Hm0Vuix2GuQFd8Q7U6n5+pfVedhTbDLcLXKvptJQQBwoclU6OBzuYltVu+p
9Ft0SHZjffovs3cJaw8GLNylYClnHPbHAobBZ0atRhPPMGH9JOYpj+bd9bKV+Cb6STAU1fM5XMcM
L+b3RdCDeehNexEcCeOs6f0tE2H4IAgJuHjDvU42JY2guk6DjgI+/hmB8WZcbZ3M8XH4j4AxxhXH
7Bflg6jjToz71KD4iHz2uEMC5iEau7kZdLattoQPlPxO9/swYfP1aJ+1WkMKDidRwrDeFgmy6+QY
jS7hRj+YYaZHCagzENunvRAubUixPjcUWy6dG4quJhf0+D8Gh16TCrq6IDMdw0p+jbxfDWhYZLxy
Fu8/7pHCKj+wvCk/nmxC7KP2YVTNdJD6gjvYNQPc+ZtCtKvm1ja2MKN9sgPpjsSlJL+3KZnHHqCa
RMCgMsJKu4T5wDdCPor2YBNH3H2v0mfiNHw0f8Q21ZHGvtJvEaNg9pnXcl0Ku+662gBurwg+ELys
zAFwyBmeamahyeAfNAFBTLVhiDh6pEu32qJQYqfr7duhD5dALBHDPjxe9i99wTdDBK3kM5TDt0Nn
TuTTXPNm/lm4AJRqbEhWmSX0u+2pBNY3eX4VaU27EXmjbxrjW4w+mw+JIt5ep5trA8PY5EA3GlUW
OXVEeC9cvSR0GjNehytTVOHTnIMrV0zSlNnRUCBlgHUFh2uV0zsrvcy5XXikv7JTkhYV1BfoGqkR
tcQO3Up6v8walI3hKrFSJKR5liS+n10LoKpaytalibPP3pL9crbXn5ucc/PWhM72OXvIb2eUAbFj
KRBtuc+TjodzqP1mEPS7RbpE1wEXTQVoXtWo72fuxGxR0Bla7uaYk6PPncaoUVJVnOYae41u9pW7
U61ePCvDC+olWFHIts5IfaqxrXXzcC8LFT2W7U6vRDUcshP02igWdufhM5COVeuT78UvD/q6DvkG
RKqYHEOw805hnbPFv0grAznfG5jjp+nLgBX0ik25p/XRvxP7FXeNHTlYt5Df5nMkG9Pt+Qvj1Hcy
OwO3qEsUsHnIwMDSFYq+hcUOyks60L2daznDjNCWpwrgmCHhD+JjQJUZIJSgbwzfbA/JBTKGe6zG
yESOEsQyeOwnZGieJXJS/j5HaZNdj3VNdo5hRvmYH6gnJ83RiZuKlAJQXvgnhajzBVAeDWF+b4xq
ScaPxKHQqgDqYqbm/IaRa1Av7hl0t3XkzI0JB1TsyOTss67DJZlCbJucJ20DRcfgLUzbaeMg4sRz
q4H1W1U2yYrGSwTZVcYvKH8Vj+NsV4TaqIxHe1ajz2xVBLIdIcKjEZdDloby0e8+ZZwYPjt55bdD
U6HmcAnLfnJA8ZcxaQ8ydHLSHryCIvLUJ+2VEgXncMgpnKjpWBRNZcBkV438+N4AREAk+gpwhJgZ
x/w/gDdv+QX+cer0cWeNst0MksTEBCRKGqHwQBeLO9D6ktS2V4loUgTIYfJrWp+VO+LH2LnVgx8K
JAJ2NhhOdj5xgIoBPSpBoCdhGejusqeoRlliztsYeCE4otbZlyb9VDestPtOeSYdAu5lb5MPlla9
5VEhzUsu19+syxIblFpgYFdFJZdy4ffPrggAoka4VCZbQ7IuP425751jh27LILIwBLjpliFRAZNE
2ZpZtiYHz3To3Q6/ABVNgC12+2/YNJlDUfnEezWxOlSk/a931y9LmcwaI0DoHwKVtxtP21jIeYLn
rjWIFbSyrLjPL96wOh0SlqmW9Hw0UHxOuzOPNwZYwtCz1r8ib4srSN8OtGsYf2ypkZz+TJkH8KYV
UGJKpgFxKX09VSBB0x0IRcLmoy50NQog3zFF5m+D52NQsanI89Ibso21raygW7dfZ6+YqR/DL9Jv
2OdGFWE3K1KtYu0FD4SLLNg1AsRYn1OuGevX98Lhs5SP6m3CnfXipSLw67EOTHnzgnnPzv88m7R2
LwUBNaMvudolbyiM+xMsqg7UIiJMFc4WTKZRyTsVKR4iFlRoYM+AA1X7+AsnCJW2C0zSglw0y+/n
5gwNSRyAi4v4fcMQ5C8e2hgsEisFptCWFQUE8hQM9Y+tnwxfvkvz/14d52v+pIPUqUV/niVzrWHH
jDpkg19sczripVM8WuznWCr9G+bLjGNnKO0/eB/aGB9nIwPeVW1+dj3+/ayFrkKPAHMAk9ZkpoCw
f/fMawfUrIhxkpn6GFCnL0h4mkps4nOD6H0jIpjYjEsj3vtpB2g6ZyLqyiQiPQ/pJt+23c5hyhBf
QOe6RYIrQp0sr3giaOKNy2Ey5tu4ljnT1sb6vVi2gnNiHn2N87Oay3Wc+4kNu+TLIaoGeNtqeYUd
f4W4QJJA+QJQbtQS9BhGBWOCVP67JomeBzr2kaHciZt0Bqzb/bDNMTfrBooj/5mR+nYE17hiagEH
zNIa40Ev4TVUViyHo+TmepfM5KGJZ4cftp4Ye2oj4O7t8uxOz8Bj3wPcsIZtjzYZOxySA+WvdBnv
48Vs76FLZmjLf0wRvrSEkPnZClLDWnlhrBPnbHEM0jZf77+a2V7xe+qWzWXM8JDUytUVnlMchG8J
Y3IYuY7qbqh15WHX25WlwU+wN0BqlGrIM+E8BqGnKZpm3hZY1cF02tCGRgYUAIZyY4LPSZp1tRCg
GRjgvJFuNaLe9PLpMFpDDSn2/8ZEZVmo6/FPSsivgJxottp5Rh7/9dAeV+zszzFteqPfINZxlLme
QQDtxcV6BTxJT28ThJaFnBKI9Nu4xRz0Yg9/dO/EZJCu6EIzZTzZGcufX++9AsKWX47oV5jatS8w
J6IGW2O9r09csnhGpeL9WV5Iz6zgROizSXHw4q98LvUdOImCp/je1HIOOIBGbQLgEG/k7lR0c0Z7
JK3LJigHSF3H48SuE5hGy4BOiG9X1XsLIDzySCWKrPWPLOe1jWzgccwm/ZyqhgnLw0ljJkFRWctv
QJJT0zY6cncW7koIeB2d/jlMvpbBFFfBJ/6CCb+IxL8/zI8TX4juCGhs98RKcN7cBEp1m4F2DQA0
vtjEc+QI3pbQLs6ow76RDMKGDe+M2a0340LMofeDsibb2ZCDp0CmJjwQYnNYqCq4Q89/6351Wmb5
bY4Er5JtmktjT3njmteD1blL9PA6nibADXAz5ti1ixhG4ogaPdDkFqUJi26pRVbu7fkUgC+P0GEO
XEmpsSxk8tbr1cyU6AvY5SsziCXXWXE6IW77G2nc68TcjF3z/FLVWJ9U7d4CpzMFDq7Uv7YLE6E1
TjuPlBO025Ldz7u4xGJIIQzLpD0l4MtZ6QOipja2/vrUbRSRtASWuMpB6eIfI63flnK0fy1MtxnJ
pKFwUJ9cZzOgBxP5/d56J0A5ev+rdmqfcDMcAb4x5ur0ugkC5Qm9fe/tXeR1+p3q6QF4N//84Kiy
URdBkfaCWyXqTBalW/Uvs7gEgm0T4Mbvy2qa32AHtLyFsr7YvbTG1Up9SwQcrAA6fbb4oFN3xY0g
bzemz5hH2jguNDv3GSmxRSCOwur4Wntsd4fK+DFc3IwQnAKu6HNji02XgipvoWpZfcaqCge1oRbQ
+bCRcG2vV7UUDeRFvoLAh8KVYLufB9CGWqa0/OKhI95oVMUTeLnJAjjKE501aAuPXxIgyFN5W/uw
I5nX9bFqgB2FFBijfXYSNT6pNgorBXYndDZHxKb+3jaAeHADRqoeUZgKA0waszgqKrH+GDo61T49
umCxfCuAg4oogy9mi2AHmYz25phhnNEKbgVxvfzzSbZa8vrRXxrn3iIl2c0Ra3M+NQOyncN1hN+h
fMfU988e7XeJDC1PD09vrJtrO03DpnuDesW2EXFXinyvHELc/tBu+MoGTa8IT0MtKpSCZax4SSDc
FDDII21GUHPtVRfNxamT21JDQv8jbDpTAIFppnEi3PSNpuqkcXGLnWkjl6/aKsoGurguKRSF4MAw
FApZjWA5tCX1fM+yRt0tgF9x5Wa6vAEkt1y2Zbxv4zNE2uySotwwriA3rHnd4RuVVr99yx6aN2i+
S1/CjCB2mm2CUT+Tc6eRj7TD/edhoiBJYv6BYlwTHPhaHvXo1a63qTfx6YYOoCgg2oDFUc4fR8q4
oT/GXQEnxr/okD79BzFHtcfS44/VWqQx4cx0zIMT+V1L/RvcS6dOF6GEYQCPbYORZz6nXicCqEpS
lGkQGc365qOOd2BucNP4VMLg5AW9irtUtYAuPSMhuyftvu7vG8fgkb/rqbUiBD9/YtX+nLB3LWKF
vNJCuPE0/kdHgrmmbjxh/jye/VH/X0fZNPd9UksYQ+IffuuPTqd/PXvfHPOYQfl5khSha9fp0K4v
GLqcjLbiVJkTkROv2lyRKeP7mOBQGfCR2Lc7ymolykBXfFszH6R4V1AoB01Qtv15QD7IinJPT8Kc
Uoc88B+Og9Bfuc6Wc+Z80UiKQE9BYsdAxgpBZ2gbHmP+sYi9/aNzZXfRapV1GzMD8u4idCftpD8o
rbGg4kniIxeyOEUwdEuiS4mV7je96Uv9wrqo0WBl1+dozZvR1wWxAj5y5vwTUmG/7Es656DtELbS
9ADuJg8pdyDNWnvvKwU7gXfyE/ee0GXW0r2pA4k3FzR+aY1pqwiCfDBGXek6c8464vBI1LxXh9Y5
e3cTxdLlU2nXxZgRq/aOhdzzArVvq6MP7UG/vRumqzPhp0xO/maP4Ees7+4m8Dr3TNzmswo3XLsn
qfKF/NKST7sqkwlWMjrsCjmaAEoVRiIlvo5oAmJFBmeh8cDQEaprZ+RpOW+nB6Y3MNQiJXDH437y
mGj9+x17cQymnQSZ2YCZ7EqwidRR9EMLLVbpGaR0xpwPu7UwxF85/5qtV3xdx69cRYhJRhvuxo3K
BmQHQpQNI2j5RW4GqO/jjkNZCqsVOPioJ4sX/rgeO+5gdaOf2ETSFZEmdu+QmGKvDgy6ivFUEp46
T0ZishQYknJ3xqdUmamrmWg3DJvDAqUt5KzNpQuo/+dBRYS6dMDC1m0IBGrmqQbbx/ydf3stXyqp
N/CvCgk+4O9KHW+JBT3H+YhJOOl4li77o/cF4Kz1bM72V9etSN6XWX+r414F66wfQju15lI+ZQZB
ajwCYucMEMFEkDQAFIvMHc5qghYnskY/4hT6okxYzTWcPykuQ+aiY+HcGMAL70zbIRyT3b69vHvZ
QkVpB2a5QIMSNpfG/nhzul45UadSWE8+rz/W3Qyr/rGH7YwUPDiUuIP0dCpHs5kVQyqAhiF9nSzd
8VQ2181eF/MZTTubmb/WImXhm5ybwL6hfaBhfT2dEkkTkxh48IZ2rcxzfp21kw4OJzqS9yWJ3b7z
s+VqR0z069PWqKEts9yN6DoSeWjscYrNpatTmtyAFRht6Q9ofGK/ph3D8xdHi4PK8iMJOazrfyYM
FXCl2BFpoYwp7RDQzwjRy3PxI6JaW21563UM3mv6cDKguE6kEKpyz53AYYe5EvjSl/10/htk6rNz
rzSSsyNO50XbFVoWBUlwvhOJfwulgROKVt4beIVZAYooXz6UMtugbV1FAZrcxXPAi46ebC8cysxF
HlMc8hrss5T2dUJ1uGbSD+FSopLioJ4Vm1RcdlGDPNdCHMbAtpwUaQQIWm27OPfPtP8CzpewNyqW
6vifALxKtykFuiZjzgGlfdqEpqbi7buWaXaw7jcI7IcJe91YtwSyDs3eKTR9yB9OY5WJtKL2nVxm
kXG0O4JITSHcfQlLwfxjRxXb4Hk6gYuo2TKPXinQaaqnMiB7g7eWBvOIYc7QB+h1/Jrs3RBX5R2A
CZA1raiQqlnlWEDzFlMUioc2cUhJeRkNvZrE4BgPuPIdFa2v2QHxumpS2lMPIc+szaLnlp6nTnF9
rYtYJ/a+2FdW5YUog8WT6KzPXOAMguWSQFHNXBat5N650z15Uy4puLwanehw2mh6F2keW5cXjTgb
9tZI3X23+im1K2f+pX6zXxT1MoBXVra+PMutP7eJ4MmYm1RcZX4axkwxNT+JZ3fj1Hxmh1jKsw+0
gP+CrAWb7qvgAHp6DPmz66qXGSWNe08F7R6gyL9g3sP9lNVeV7stZtZiSCaeDMnYTcfAKDELW+TZ
BBrczTfv1quhRU+bDt551FgNGsGG227bDiXfZEhYFb2tJ7f1WOJmf9n0Zwpwtq3etGKF6sq/3KJn
k1TzVcVbPpW2xduK/8IddCce3mAI/4/PCbFHqTiE/FRGcA9l92+VkmYe59yoTVObGanny6q9TPbB
xJjJFF09849a/1CKSY8cTC58MXUra6k6GB+PaCnXlGTVRJFmr0C0HWd6gpr0BIfQstwm4ZJvxr/a
7IvkqQPzLQBXwLLwk7k8e7wjmdambaGUsyIX/GlTqp/a4P2nnbc00r4SN/7bxyB4WW2J7vek7gYZ
TLMNtn5IsQMHXI5hC644PjjSSZDAHulUrkshnq6RRpApmRmPVBZ5qMfXSCdqQ7/l7SPBJccFQFKB
Y/LciDKm3ntUBKJ6PNHUjxOGovtCetscXRGrV3XJbYDPZt21j37/wBq2EtuFZ9UK4R3rl3z3IUMf
DyK+E1arKSRb84ZlNS8JHZSDxr/OhXKwucVmNREpG58ZXdGZHBjo4blSDZe99y0EWmHkDCTJ+Y8P
Zi7jZCL3MCDzi+ltkIUVKeZQrGp4Obga8H4pYLgAdXtP0HRHfH40CaeJMjKQvLtfaHJhO8q5D51O
9s5WCnV4qPk9YHhEAsSa4dcASxdWpfHVEyKVhHqdvOiolsrPXE+yL/vvBssYbTqrZlPN80jKLf5m
3gLTmlYqunHwKpH8z0P2GcIuOpb52PKYo9R/bCkoS96lBoElxCBC3ZMkJuUrPWWoaR104k4LgAHb
6wN97qeuakpduf6cq8/tvG4h6MfuaHXvfXjfZ94tqH4Z91OjlgURM0mwR+Nmm+WLG9M335Ux7XE4
je9pkceUW5o+ROXZ5IDrUEtZ6KTWFOMnmA/ZrogCevLIfnfRljKDHpgYWO/gmMg/yINGgykAggnz
4A5ZOaYhqZaN5EZzvo04wvEAwABxQeWwFQMt+XUfO2C6Hz+XOfGZOuzIqekg6FBxzKNGpMQnYplo
x1zAaHMCXcCQSMwR8dpqovID9vnwhVrwVrOTmbMNdn/H7MRXdJcYGeMuXSQKBFcSwgyBpwL3VepH
WMt48z76+76JKMbhoBm65i4WlaXFMmlyVdugQgx/r6xIyp1WL28O/5gAwyO7vSuoLgOb2TJpZLX2
jh0msdn2RMtf7gjySAyK2foALSkOWGRU8TK9PCYxtN/5WEdPHzT4Ah2twqSGE+eciziKk0JIixLu
uwzg3MGc5/Cr45NAbKh0jN71sYHdWsHedm+bN4VWvoUyjlI7PAHqb0CFZDz39kbk0LG58G1MIUsq
TWVgmDRTS989YPtIONVMiXWRGmmWFaHLqIuaZdi2dBnJoPemgKY7IU0OACB8rr2MOitxuIvMU7K9
7AewjVEB1sKVy2Ct/USYSxp9KYUDRW4TR//SbW+BL4uPdQo7y54c7w0XiwJxFhKpS2UZ4eImtYyE
qMLFXa75vzKppdJ24eu2C6yBYgfdqtIDfMhTnSlPVyOKNxMKhvEWg2m8mjYWf6elj1HjUBOSA6yZ
1x0b9UyBK4EdnJPqPNo3VCT5HRrgsKcD1NUlflc+dB1wXRlW01+h9qPppydURPxyPEn403VUxn07
D1HbnJXN9IBOsq+g77u/SDq0vyC+0uCCBReAcbNeS++OeV0gFvh/ZBhSnFRUhmsxR/d0jNDinDZO
ELmvBQBhY3K8fJ9jod8lpciU0X+2RYnkq5uUWXs3BggRgbZVi50CKQzDXD5xmXr6LDLZTrv/N/WK
2PH5+Pepu1glCQW5l6gheLv9JdGtndAuVgvP7eD1gBcaN6WPwae1JSJyCJaY5cADXACrInjJL8d9
GQ9tVay+g5OoimurCx/IoGVleTNHmHHRxcH+InsgR+f+a6egPNrHTTHVFWoQ1pxSI32/xddg4lzK
4LWxWVmlhT/L4rx6rqjFEHmc5J8ttHhtPEIS92+NNOr5UOPWZgBRk703Plp39ucNZOHWiztUofes
QuLILJ2tZ0UCD+4+6WmTsFC78So8CFVebzq1JuvZ3mpS3wQwenh1LDwVah71t8vskWndV3MQoy2J
31r788VwfkbC1TqGEiXuA3tWjdx3ws9IUY67S3EoEBiaoKfWZ3syCnZcvfyce/JjYisKQaAU5Vh+
6LyEGA7QBy4+kRPKlKjxExxfp7DprlwvnXtsaI80shdQWZzrvoWwlwC1bM7BkI1+dN3POMu5Yefb
hnG2Ar/G1oXZ0zd11r9G4phWzqqVryJyVvHWlXKKNwXkaeZRC7l9cBW0u9M1rR3zK9vsaO1mbaNz
oT51XnCDPM06WW6OK4GKfS1RGnV1CUZynMqZytgLI+OHlV74SypHI6dtUmwtEzSMntXJrplF1T5i
CY1ePyWtGC0yiNuR2b0RGHbztqsoxkLM4bXiIeKCgAhZC/aXxpdkW4+YYxhtKxtcE32a4vb4/Ncu
KGlVHYBA4Nbhw61XjorZf8BnO4uwhJkYNROUB5xkFA1CtPi44otGpu4DsTQkEKPWOZEKlyeKYCDf
Ncadn6K0dHWCWoT+uJI0NzhSYwBcJDksZ05fjYj+crhxnIt1TSatBOlCnshpABbkKGUCHWZH1Pki
xKIzomhaCEHQLudWG/mI6/en4corviZhXvExvD6GWkXdwW1X13wvoM71eA02zJm8TifEJP+nIhqH
dUDnbi4wpNqm4uvU6L4ldIuIp/PWz6/q8voqVWFysfl/WsvAIR4pZqM7Ri+CwIEBkyCuHbKlTb+s
Ocbn0cNwioH4W01SboY1xX1tqfz5bEQksdB7a6BOUaOuLaoeOWB5OT/ichiGy5ZvEzVUT2NgtHh9
/C0yibSE0g5BKXLQoF/DliWxunp0aLushrZKfhmEyL4QqskxxCMiW1JMqhI4FzxMigTYmm0MU9ey
r2siIQVB9lNPjBSkfy73bg8NgWvG5Cl2yEh72J/rq+HEdaxGJz3fEQJ6oTZY2hofoAvV/y3WEzXv
GE/ftxLWFWQDAWjz6qsVaVcuNZ1ejkxiUk1VLas/cW5xtNdUunzNFwOIOMIJsKYhI9fv6uOPxMwx
cFTvHwgWEb1P9PBQe6dnrqaOhAG+HZQOYxZuGiaD9Iiry8uGsxd8SxrYpaKLhwT7juV8Vzd402u8
ZZDvOKUqw0uuDrPc3ywh4HHwydHWUJN/WBuTtwkC45xfaswibhitPAveiFIgrRpUib3maw+bvnsb
nAGfPu+IoKmXhDWzXYa1S42CyEBjrWIlrB7FDguKJz6PzKttUgGnkKIWNA28aZtUx+4JWxHG2Wis
k9TMJAofV58B+r2m0E/AI7Vdd7ttKvya3EchXoRmwryTtm1ROaCsqj08FmTQI3ye+ajeM/Oj1pZR
Jy/i+ZyJ2WW6vS02t/XgMkcGVB0KvyNakW1goFEMROtsL6kNis/s0zgwrpRvPjEB9Baj5jf2FPWc
DFChFiN5840m5xKTyZ7Noem/Ad8n3f03SZCnvs5uyYPKgazpLdXmguIe9oAelV5xsiPxpC/Cw476
Z6JXglryL01DITRZ8ExcDoYnk31lVG4c3PMMOfRFV2yl8t3gWEBD2pd9YUcgRYV2bnmEeOsA+EdI
D0Tvotnljb3qBChPMd5yLl3yGykZa/k+cMPwq5QS+mxVzG4cQthRfIndr5ciTpCJC/d04D00JyL0
1kce/Rq6j3YU2EGFgRwDvLDxUZ+s23DpdRWXej3c2fWDh5KvGrslMgyHR2wnN6t4qPnYlgwGHII5
h+zJRmYmoweSIFFVriEw0+o5iynZJlb1uz7l+qXUndzOL4PlS4wAP4XobdXTQBNz8bmNxeElyjZu
+cN4ZUe+Mvb3navknLkJZY2EEJg4H8Dg7LZZx5LM9F/FOw8qsCXbJlfpUoK9F/TEwBQ7Bvj9hncp
Z6X+jwrYL4VCXW5ICxv95cyzcXr+E5TPbc9bCBq6nuC5+FEuTtjbPHBxdDIMisGsjQpKGUk7VBjF
mYJ6japzu4vph4pKYwJRo2zSBVZIB05f0SRuACeCwKFyRhKHHJRBmGXQuJSZG8F3NVV/CBSnOZXs
4OcgatEFPYJNxVN2cTpPSWD2EBy9PMA6nA2OkKw2u3J5oFJr2qc9Fl9opLUNVBbIuQj7zyi+YfW8
SPmoFUZK7VqhOEEsNBB2c5EKK2mhBIR6EqrSbzSd50fKmYFMzIy5xW4DOAfGIS6utp/MJte1v3lG
KFTHECRe3NK/WgJZHTV1K4SFpNgy/lnE/AHqaj0evTCHE3nVI/4fUs7YkiIdQW6vgViExdqMPA8C
irnO3py9kXL9WOYzbAzm6ykm7pDz1U3DzO3w+7rpp5lAkYcrhikBvJwRJ4lS84uK+nnxqBtBMkMu
R/V2/V/0ro26pogqz1r+MpNH6AFP9LEyYY52CoqecQSKHkRZGOxdjB4b0diugsJBG51xWPtZQQ2U
vrMJhmntDQTzse57EGECdZBG/SYMed+Wh3ykHnUwbnUukOEXD3VD6TBgVO1uyDtbomE8zodshicL
vaoMpH29YFj50VxXTvW3W0MfdfFNog1Bb8v8XOWQiR7t5xdMWIJyWb8hiCeMwe+rWA1CDV8w+gPA
TR9hAcOrA8jz67N3GAFtA6zzK3GxhSaRkVY//V+k1tds5G43+xMy8fbUvoigNQJc9PSPjWZtKGVn
LkZZnBOVCiHQkT4E20Cx5Y2fXMJxrQ+ZizXoHjHAWcn3sN4Xp4kJkP0EJ5yrN7k9r4CFcxGcOoMm
fHqYZD7f9YKr65XbzSs7cQ/IzbFA++JZCEvngmwSyPrMNh2eirUpyrXCPWyF9BR6Iue/KM+TzlgG
zwgmONKivsHGAtUt5EJJ18OIDXLKuvXfXEBUHY7TOqbwUFBgatj8uyU9ItB6tr0S7Wsk39Aa20pP
RuX6TLo+SGxmcT7gozH1RyG1wt9bajLY7pOEjazYkdtNVvJaP4dWuVZJLNHhVpVr7cSMmkVWBJbE
vmJl7XvdO7oqbEhBRcOwBK30BisPh4U3V17j7SvnMNUeYxeZHaJ48FI8NimqoD5bILxQzQ33e1gP
NMbB736LBcfz7ABOrHU+iVa1l36EZLN8FaE85FuE8svFJMnqSc/e7T4YduU+fK6+seC0Iz3liiED
JEF4LJOFfmQWHUj82YyynEfdGJAWo+z2Mc9PQSg2Lyq6jMtMqVXN+tdP7vTuc00wycrwqD4FJpcI
OI/ZgDjKFCy9489CMENcxEslxFlfYLlBvuiVCTnfM0+z9ExYqO07FCpZTLlD8d6zNyDiDZ26EV4T
iukdRJPaqV1zp9PoaLwCeBMjIiuU9fcZp2zer1C9APrs8SGlUchKn1MJ4K74J5YtfFyNzokdzPxV
iQ6xcITVqeUt6GoC1HNDVl6wZyepg5CIcXO2hsc3t4h4SiZiNY1GNyFC3p2Ev5mwovrtjXwDtGYn
FSRIg3Po8YIqeWt2wLMz7pyLqb/tmuvu5xsUgjkcvVFXeinYnbIFESPPyosyEVAAuntqZ3OOaxeC
G6hLCKVeNKYUEqVXpgeKU/luZx7c0hBbKdgjr7tfVkIeEy42Lsb7yth7iX5Y0e/6h8ydygRUc39A
06jVUysh1MxQVFS+fyAfwMEy9zPNzGmXYkj+lx6Yf+9EXCHT0jjyGfJyTBIhFCXLYH8B+co/YCt0
aX+4S5VPJSOfVmJwIF2WoRxRRDYfMd+UK+hOaQpKDdn4QGSYXJNCsZl5ZWoo8bOsSnVbFUpE4Z6N
yICRpiZ6g1Pn82gbpGTt4viQPxrTQf0ZuVnJ4fN/D7ohG7hYLPYkS4OkjQrgPG7ffkvkSvMbh6KN
5QnROJp5bf+i0PWIhLxbyD0ISx6PNu9k0qrT/a5DKZwed3b8ANXL/fd2exJDdvBX+jxjwOaPUJLa
lbD+RC1RweDIyPbxDNKZxZ1NVamgk4Xv90oAF3GwZT92FFnDyxT5owIBL7R7PlN0RHr31ApEB4dw
T3gfUFd5Wu8wU4/vBL8T10hHtPmTLU4JG/g9wpEqBkXgWrVuvlpxS5ae90sVcW4iAO99w8R7J0Fb
NkOM4mSEwo2ojrvLJrSFVRgQYujgNAyOgWu18nv6c9BGCBhB0b5JGjwDvTtN9dZBYLRzkHVVe/4T
RRK0yiyABZZeypikMTwHQfpxGQThu81s8RpHaE1Hub8acsrK8xvVvu4KWsotUSjkFZGzXYgi/Hbv
aUDHo8DyCRCqRRzL2XuKSj/3uvEfOqL0c8a9I71ROi8RcDRi0fjgDy84NYSHQQyEAzPbbw8vT7W4
FmY5pE6Q5qdwNdkmXbceQRHC+qI16Pay36hQGlE8FVxCOqiZ5xx6NjpY/ggTn9ThcBvqtyRiNgTw
PDWbN1PFw4xjrKTWilX6nJH3uEuBt5AS8zE2L3UCqU42oXFM+EwCWffuHHklkAqzPdn7yH5OaFUF
iH5giUnoUR+WjTDsBZ9+f9CGchDPsKzXeOcQM3RzVfhcVl80qtKshEmfhQW7OXocSRYkZ5aUk5Ky
yjiI2gJUT3fL5DKLfkVKJHDaPTXSdo4ZltKfttduGC4fh35SRd7RtNuG/Klc1g+Zy9mgQhxJ70HE
ggg692c4jr8k17rpLg6iv7wXhENM1Uvx+R4apsxX7L//CMbQg6auxtXsSe41s7wwxUWNArMgl+IH
2h8hlayy4eB/r6/HkZzln6UwT8fK5ZkJyfFsX0w7R1EE1s8g8ICj/vrxXOBcshxJ/rxvhxbds84r
b/WXm73S6+8FiXREu0Lw3fhvvxgk85mNxfSmH6ePkJo13t9b8aLiXWW8jc4amvIvJLTURIuG37sp
B/N1iUslB1AJcp0mMZjr/HwzJdAImAJ4ur6WkrKzJQVlT3XdRm59YDjOX3N1Wbq80m+zBQjx3PY1
NxT+FtFRypL1oiYK5DSbb3oNVO4Sd+Du1IxTwZOsw5Lph0/nmXTR1roR336mRYpz17YFpOSvf/w1
WHDQZNtBPfn64b8EhsUbhXkLHpYmPRg85pxTMl92qPvO5Rkkvjk6Uma1yfqMbFL2dvlPPHJeciEY
iJeIFDHG0pIPpLN//dySNm+RrzcZah7xnYGBDtJf8pn/eUZ8ACa7iAqOQLMUJG6t+z1mAih50wI1
VebHl3XN21zzP5gDI9Kz45igDGNjxGVU59JI4bOC7bqBzXNeUVWNgszeFnvJzHNu+7C2YnHEX2dT
6p3D0Qq/7ftw4xqJkllZoGWcXTHO0uIf8AgKvsRVZK42c2OmSstdsJYVpwpOWH2cygSXJGjjsgW+
GKm9KXCLJ8KfDaI3Yt6op+kcFp/s0BR2fo4spwuawHn2ISfQ2AA/6dPPw4tFZTNhS8UM5Qw3+Tie
TRGL4verD0Cuqw3Q8JtSPvZHFjehwoSAv/TSZt/c1KDtTguSTRaG8o/Nx3eWiKsk0SD4iKRFTmT9
4FA3lx5LZpUvFVoevck8ONQoagACvsm13/KWwa/2JksfbS4rLvYlX/u8HsjDi/1oROdExQaWHMzV
Bm+uuhiIFXQoaaLtGkukpfsu8wsS/UqSqIfMB5RCvVdVM0ffGWGH76u+F3SuC43zIiodrlfYn3ju
tsrC4hFZmK8p7s3hfsW/1xsLKpWKo0e4NuaP56zi+gFd4e9lgf4y5vZrLLl8nf1BkuXw5sd9p4Pi
UjhYic4lzNjyRNQDMBu4HSjj3LfYXhpEjhXNKlWfRy6Y281QqTRQzyPQm3PEcDpgoDtnbJyWsiQJ
8KJMWV/YsYazasD2gkBgAIlhz2m76PxYA2/ZoLY3g7KOfdLbtX5LVC8lJGWz14o9bt32kjTRy/+d
5zXxGhMKt4x2tMx4ERH5olHRMUl3nPw9wrCuiYj/NBDjS45HoGJ/cflBSHcePSMEQNKChWfGyHFz
atkP7W+tdpKHqyoVTHUhyPPWv7y4kfbZS3ELraUGfWB579uwrJ+GMn9PDIcPl8zBobPVHY+dvQhM
rq9+MXdX0rcbe13kI2WoxedHdMHJaynA7Mq8tT/cEdfKYQwKuA/k8tO3ud4t270hS4UhlqKY1CRk
E9fqjsfdXNt3RU4YO6uvHpFITh/17rNgHtrdqJ8GlO1T8Vxf4aqeDkz5ImGzTK2wepBZQtS7b5O6
x3MELrspDOBQO6hCE067MKIREqY6iRrCP6lD/PHXKEwOVlSjwedLX5SLKWRK5MJ89uggubU3mGMu
ae72jB2QdsNl13AGH3fRnmxGCNoVjbwkuK19yWUgCIpIQ3+r2l71rXoRe+6uHUnlCVnmIxEU5Tdb
z1eNq+xOZ2tvGRRbAR95vjsn05eIU+GAMdH7WagA3FsiDtAh7x9vUlC2R1ffr9c/W21FAcBa3QSo
jt0GPmk2yoVXDETw1wG9YxLvSE+0MIeKSurbbY/xRi4zGIkb759rCA7JDAzAEB3q6kYULxx4IaVA
2HbY5T3BYhgNYs22S4B8v4oGzxyzDH//BGxYoZuiwt9vVbmLwnsI/l6kBHclU0fTuyrSwNHAg0rr
CTNfHPUP76OJ2Wl44gnRw2h/O9NW9z+IDwVz7JdwuWaJnZ4Q9Th2qfdvjdInwWklkvaciyU2VD0D
TnmS/M6t3QCjMS9XXuuQhzoxF6HNT5IFVV22iq4DNlXaZWEf6IzlKMn1R0YoRSEy7DeuEYcQ8lnx
Bymo0OfniDiFZFk8TAWyjSxdPf4ybIMq1Yo5ZyZHWmhM/3a9kB74ucEPDroXtPfPnfdiQU2KzrZR
leLTUY+VrliLua1N0ezkDx5wHCpQKe1YfB0956u6Hpu3dW3PKognXsqm6F0aiRRjinnWJzKYvjty
BqH3Iju1dFXsSzBBEDCbnLbF6jzBiTWIvqfjqmpHfMtbrrf0JvNtCf11k+RBesmfx0lSpUx7YDD1
6xYzz5AoFf29U0wlwZm/oj6sMcEKnS1lqtTnlqMKGw2+78jdTqDZ74lv/xEp5PdV2Th5nwnMeR4n
eD2MVWCCVe07sTnM8Ljt4smw0dcFL1mEc8pNm7rcM91wxfPwq4q4+cL8p+creVUU0lU4nSIAJKDf
G+S62JRnAhbCOme+iI2kR59lRqShnRMECgfzlU7cf9Ng7L7bxiPX2yR4bX6VJyi0M8UkSXP+gGa3
R0MKN38Vl/SOOzaZtIgrJR3Jws2FXehLMH94P/hW1+PKLrelJgCLIvmVeo5Q/wVn9vGkRk2gy5MX
r4qa+/kxWNlqBp2qoL6kpPR7VOhdm1IfzbhlUVJ2CLP96cItqu2m8OtXNbXv2rlzU2KxSkKS0G1W
/EWHUiNSZ+MNr06oXgTiHVmLHQSis2Rz2jBwEMlFEBAEY1ioFUPiXXMzZ841f6l4NNsyHpQ+llEZ
ZIBpc/jaiowzepLQLVnxMDhPFnXwHF+t0AoZRumJv55kdi/p7TpwjMOlirwbof8sp23KlLgcxN+f
3P1r5RGRB6OQRgs07Y+GVI70XBjcrtCeJMUkQ18Hf+WyyeLx0YpCdSsXHzsR2FxLfV39OgAm01Vr
xjUuqS8BKFqVek+hUUId1oCF9J4NaILzPGdZZ+L+MOIE77erN9k2zuP9VO6KN1WGDHMzKyR21vYv
Lxcr8lrA7rfYUzGsHRQeCsV+lHnLUMJBgNQUsjtn+umZAGxX1kweHEy/k3kAtnvF2YTqfOwj4kco
sNpMMKdBtFHdpYowEPSPSUuonYb0GJls9VTkW80xkmtD4E1GFFbz+rlNg3is+WJ4utt9YtmnNHua
5QeQxfTRlemILIJfL4Jrib92wtZzIyyRjOyZz/CTAN+OIYzeylNFW0VefJgXnJyxEzgX9vyusMsF
IAZmLyc3WjXuwEG1f5m8UAusdTgMjk99OioF6XplsJ+hZ2wvE4OD555Hj51FkEBzgWAJvHresFzf
QRF4YwNj53g/AiIWbl3mAH7UH75tDwAEp2DC1sOEeGjtn+W7wHRjS4bkr7PZOGESnFhPkVDcp8h5
t4kGotBeNQwPu5c2FjMDeYED/cyJWqQOdi982ROsU5E/GQ5bkMNjJ6sfXx8GLp/+sL+EQIkUShye
KJtC1waczui9VYCff/YCldW47fh5ZQr4s1vOEkOMAdoAD3mu1nh5O4S37bqWvw0UtBg3ow6GvTlp
FIIgGZGBm17YdOE/AY/pR1M0PgKzbBn2YG3DkTl1p7J16rJM/YDamYxZZciBgPSaYHBuxmHaug/A
yLn5j9f6IT/+HRBL2ks1cZQFvMrU/GJHdft84IOY9UG0xYIBJscOhdfJE9bxSk0EoBMA+yyiuFpK
vECxfhdzxzuHl4ZFHMkzVsRUsuwo4YAxxc2r53TqQqvm+fTAqcQhnpvJ7npk0V1oJwyExUSKYhBA
2LEfI8PBvtfrk2qgy8APfR2W4+CwMQt0aG6QbSHHzFXK+dX9asccSxqCmFf2hoYa5dN/Md95XVq5
IqjNnjPz5L1IIN8vtjeHfjSBJohNMXb/vYDmYPjk2dEIanqB9BmCvH2ksTcsJPIJqCJTIqitaKkN
ffPUa5WRSFj1QMzUQS1Fz48ve82GpWK3H+ZVyQX1uPfhnFMpEEUySGp2HBT2FhiU/hU4hQmvhq8O
6qXBOpJDm7+Tq6ENY6D7yOGsmKYeVl8tGojZFedUrYsXANoscmhMRExP7mQ/muqkCQAiWQNCZATc
jc2dScHWSlf6g95OQL4msF8+EXJYCX+l9CIUqM1eZ8qB/MfbrBuYbPDdVcVq9ZMvSKc9I4rTfk2D
oBD9+fsBKnNcHT7TflIL/bdDT7cJrnVvrR5Q5bFQWAyQlwiY0f5P6H1bpA3fZ7ExZfOCJMm3gEHA
MjVH2l92yBaHBFiseytDVTZP3c21D547uPkQgxFQtLlq+N3w5CyKg7/G1EZtLYj2pwc+MJ33kmlw
EFCIJDHZm7tVB4CrF4ErxMfrm/us/RUMXe9jUnH7P0kQkNlUqCAmhYbGWQxk3V13ML5RD8o97wiS
+pwIc/BJhKhXbkRbLMFjeCINCOdAezZAyWIJ3+apxMhTX28ximMLx/Dc/TwO68m4F1dETIlzcLIL
XKgWXjDBaVOheY/Cg78CmyVqEdB7DKgzDD9doUBRKKfuMNSLUt952AYiE4Jx66xipHNPorxv+15y
MOIAUqdfop/w74YSGvsgvg77J0JIrZYWB6mJB2l+RoDM0aeA0LYiflxtj8WIIDfr0TmQpS/Cd2+m
9Bf/LSLvGnM83DZ0kNEpWDWcEhF46iD2XS+fSCnVX/vDzYauixifykYxljFeMgtTJEGIvaqMsBc/
RtfmmEaRxGk0j2Nh5ESu884LpD+YpLUd1RnZAx3BBTDnt4EcTLCaW7Dj4eVLiliw/dJ6Ev84k4q2
CqRbJFc0i0OzFS7QpVVeVjz9FZXpyob98zYCj9Bo29CKU/0FIT0ZGvz0qHOB75nlc4sJw6ISydbC
K3vkRM7bdci3Yc3CYNJHSWRkQzo/ISvRvj+O9ntrsDXCcTeTw8ipYXKcY2GZFC0yAwbytHW+pvkF
xSTbY4/PCuOaf8G3CkOFdwbVF8Afnfj8wtzoP4JythuOiHA2ezV/jFxTrZ4zGuiDS27w24UlVJnj
07v7koTLsedU2H1W2QTXQVlB7NozqpEsic0Te+crxfelui0mWom6szjIUzR3QKlYbhKmHwrgSu9m
UJ6UZMOYqj64RRMGKfnJ8pGJSq2VGCukGS4cW6FRrtZVyM4DrTCYBR9zN2iYxy37vJ3WMJhVbY2X
RWEaHAzxQQ44Fe2LIUSf9IOuSArtXcngKxqgqP0hIsszUsLf8iqazDdbn2RIuBYpjmrYDpOMYz+Z
QjitYe25YBZq35xJLo1pe7F4GQa6aWZfB7DHMnM7yNIRk9c6Z4LLvRl/u9ts+rGSThpqVpmlOKGD
RS7lKcnar6SQkxfytOJBoa6SSh0Ftq6TEauuNlgiUJA3B46w2AcCjGXzCBFXttynPxoiHSxclJA3
CLeL0L3PpdI7DhbhE1TiWk5X94wI/vm4fmIjDF0khjsTqy8qsAgYo7yWGTJfCqEmS9Cvcxi/Adu9
IJ7MSuQck06zv6pC29u0oKcCXDDYMMsMnkzw0CBEYhawGziuHAsREdqk8tsSesoBF+dF6NME5vRA
yxd2YT59/vc2foVD4uq6wUE2bgUoNk5y6TapGacmT3pzlKqZovR9qjhRp/66EC5qnouBDLUzNWdY
zWONmnQ2RhqScAtCZqYSYtJXi+umJs30gvKyOsMyU3JD/4CuQqzL4uSmacdfitpSA132OH8z3pmR
Gor1CNcBJJkE9HmqwuMwW6X6fbUW3RlkNK39cuO7FNErlj/hGEwT51ub8CKgtAvbcGWRkKxIc/iz
hQByUUq9ieQ+efaoaPOTcGHBljpCpm7jrhe68393KWuUCRKjNhKcQO7GGhgD7uQBhlMHDiJC4Jmo
OdR00vKEq9c3d8v/jaZGqPQCvZT94oJoXrnNMxBfyb9wtLIU0rFv+5yc02shcxxqvvDx70Q0X4ee
ONifDuzuq31nhwc/3v0uuAz7UZQWTVzaBebgyJieswNpb6KmhFjpvWfhGERYbiPmUFCWaHWT9vfk
QHql2oFjRxODOM1Nyvy+E3AIhu1JiMef59TldJlMlJngrR7l6RGP9smcjMFe+eiMGG0EX9Z56tuS
NyoEHMfz8gaz+wM4Oxj96ZWPtAzJHB5jAoAM35IJARYuovfQRTZx4fHtlea7dECp9mQXqrshmHBS
ei8SffA3Hte85Yws8Kojo8IwNtJa2gX+GI2mpLtsZ9QrjQO1fssh2N8fjfznVkNJyq/GlFOwmg6Q
6DXlLQ/K5TRS8ubcO7Ye3PA4Z2fgmzTSfjOi9EvGDPDoVrPkOuCKOWEvIIpnroIQ/g8Jv+JDEhqx
T/hsBsmxTOSXHuSHM0FPH4LVyrlunMT3hM3qs5ohlJRGymTORad7WVcG9d6HQ5nRXJ796VpuFSbn
eJc7RD7xMqkwfW0qABRe5CgpxtozW/Pvc8L0fQ1UbhwKeyLz2osPaKG+TFXtoWnZjlpBp0+m5VJ2
UIrBm3phhwVNipvOqiN97Vc9a1R4ODH4gU1nH8T4bAJpSIlE3KpqkkdAsW36xEpVNm8yvF2Se6rc
217CWAsIRaANzyGzImgvP1ty+hkgHEMmir0Lp+792u7NOwzdJ+o2+vO3lb5E77jRdtBYrIqLglmH
n5hFHb6P5TevOD7IAGbgYanfMMll16mlK6I2SMnEODcIg/qN19DdkzienFDcpZ1Bsph1ryjei/e9
Pos1WfKWd1RgOi0ZnvVDcyRdPtEicRmASPdgt5FrU55XahNiecwCteou0b5Z4plZiqQq7BOwJo8G
D1h2PbcTTovzFmCJNrO4ttk61zDFxRiH6E1xhJpeo75kcy21TAv8xJ48QPQo+1Je6+OQA0l84ybx
uxvbB2HeivwNvF2CNje8OpfjFCKyxwk/dcJj3ln2mAyaZ0Mpm1Ga8G6oMMU17QzxPUVm4k12TbPm
EnbZ3GODpvkPPX1b/H7Ub3wnEs1KG35TpaPetk7c/dnPBWZ2BuxIkcWRTE2daDNiSvjlBmSpsdfz
nb0h8SYDcvmtygEd8Y694JeHpoLJQrMPwM/2MjaJgDSQ2fpz98nesQIBF/YCYrtYJDCfcJxZsAzd
6ApYtWZCqJSwqvmVAkC3OeOWjTm7Pcheixo3GPaMtEr23mIcPQrSrO9v18AtNF+9q5KjldyThCgh
gs9bUaElonbwPPkI19qahkufyzQMQzQIjO9LMsRqpvzq4M0371WD31AhlgTIFQfXIDl8tPimqysZ
6HQRiMWQLXwdI6XipQ7NL8MdkDPel7mi/en25hWxUZMXz/ZoSHS7nPAbEtvNOqerbGNmwxucZNu1
KgTvBe3IQxUwcnQgiZ3HLKENfaONhUAruXrFdJ/GJuCwLp687Ju7XZGnrxAIXBORHK0dWuIl3Jb0
7+m1B/POgBzID3a0q4H5dfPPVAl1lQO0DmjraJ4uoagFiP2OTyZWkqCAKX728bdp/ip6PnvbKVSx
6XNHjFFNXZxfMGy1NH/+YBEJ76RBLUWYRC+/4djl24GyNJ+EOwGkILMjGFfGlEH7QIzBsh9Uf0vp
Szl3p6jrtmr/o5V/Ued9M+n8XPU9xpjcDertV7N+VDTHnlaDS48vg5gI4QXBIde/JSJLL4MBg1eh
4x20J5nnE7jyV7D5EnmHXl3Qax2A+JTTMgbgdC3vZHyfqg2t9KUUhGpL/gReQ4AFthtjBkoGtGfq
tt6dqvNPg79KWolsAKIbKAr3M93u6N8yNENIkgT6ww1od+3Fk2QoagnnJ3y3HlX1xNDfhZZ57QMH
rGfOk8wrgiMidpGyAXaD/KLADoU/UUSr9rcdA2pq8XkMLNHQ1Ft6bwqRXnlqdJ67TTMtwtHiCRFB
+ylp/IV1Or7ZQ8QmB9ct0JtRIskrgGTzhW4XAcN8f/snFTqhI3NMPp/3aaJIInsWPLM5X8VMhJrS
duCghBR6N/bGipvhjUGfO4qx9UYlfuNo1R0P+SygCf2ghLQE1gSNMq1HRnYLNfEmy79oHZpfncGo
YtzSDxxBASjH/9WZ/Qw54RK0Lb2mKdC8ewXkJpeumVVzwwGljy2yvQp5L1Zi3vTrnmhSJNJa8dBo
sycWX5G2p9SQ5I5rSKTrgqmG2Ej7lGLFXZWGCT40lftnrzSXucO5/OjWqQfmRfn/rOe/9dZpzmyc
1OubJfLbzb7UjkVV4bK41vpNjSPOcdzoeQhhuYMpuS63ingOAyqzPrmqZxA4yXWKZzpeU48Mqm4h
YuCywfJYSkDDtyi7P5wyhaal7BCCJEfT0HSNjp8fVGZGVdE35hv2c9tl9Wl0mL8Og+RWe1pyHQjh
oSBd0TRDnhF6S9K7KXsVcjp8qAAwOhR10s/tOcdcfyueMQycgwLehEBV38IWq+8qrFeZqHtiq+uH
8uQOwigIWBv7Nz6B0vaMW/NxeyXTbIeJKdcPsJLOJdjWE7KkF+JXfmIJGqsGkNJ/Z9VT51ZUw9RO
+ItlFQ7lk7Nc9JomkfmIlgN6tAOUda4SysheO8LuuWVLWuxgcOEgs+t1at65IuUwz+EOncg3Nn/q
ATl6KabMyzH7NEt8KQqcV+Xrlj1Nqkhu0olNR3ErtDgXLLDGShBV93xAOyIZWxBuNilUC/Gww/bN
RA/vSZLDJ/jxhPwcYhSE2uurrulOC2ef9w/It2x0hGm+Bo9jdZD/4LE1POxyxD8rJvStIxjOPx13
5m+4uki1G0OklrHFdPqsdVZ5Kd2pahTe1r26DRBi09p2iFsuqPzKAtJLqxhFaoO4DkcofitDl1RX
FME3Vk0m60Xap+EZ9dZ6y4x0BQZ9Ehgepovb5/ugWFV5VNuR4vutBrXUM5QGbrwusOpJg9dzE45r
NF4RgmcgIBRpx6e/p24riTclIQ9kxWoAqhKXPGxHzC6B7gDE+pGXLSS0gjZ5D0pHDaqSgrSDjfos
EPqmqQKH7lbKx5vvrY6eSs9aH0vXSDUFqdIlfljsi5OSu9L29NhU/VOzkmi9FZ+g5CDKU327QXwD
mchH65poUb8xDGofF4i61f1eG9M/Druh3YtCSYrqbJkwf2SlQ9mcIbVfmlkvkM6z8ybSrqdnoMdJ
D+n+hZu7rlfyxq0Y/Sv+MCQQzZ5EzO9DB5UbteeZcm04xjRT271NNy0Y/exzfHQc/h8Z1l1RYMPg
naqSMZQtBwfUKSCsOFWO3NOH/oPaA+lj5IoNRotf8QTOcrnop+DhhdzNHpCSf3cTvjNTO7ixbXZM
HLVWxZlqV2ao5DdCdXc6OWm6sWsMjyJ4XZ5Pdjr80t9/8iOOdaTpTkmcVe++pSM47BdbmIpyUYWZ
jfOUpP1jB87Ko7ifowFoYCERQQ5HtQhW4Fyze1OydjNrQLEmW4Ko25aC4VawHt3I9nwqde4C/cBb
2DGEBTV8vfCXo5ZZrg5YXtS697dFTl2iVcYhIosVsii80z1OomBIvVHq2YPxp9Ox2eUQq8tx8gcy
/IIzvshng+5N5LoKbpkfHxKOJQ7mUJSUhx0s/1r9fvOiHk3c8XwRc4TpDQKGULIbaMxWeqhcKB0u
4ErOQos+J7ObSYCo3vJlrDsDwMBBfEM2Brx1ckcI74LXj5vCA9w1f5ny8wX6kz6DUotgcceRbf/r
GwGUKcW6FGacWl5O1pTxA89rBPNBSn6GA0joXE/6KcHj12WXBpMaSTIWYYBETe3SgBBoY6UyYh6S
XeFzpUo82RrvIfETCizyaw6/OdoI7xu0xXWoymkxr14sPD8750Muj37P+1UbJu6hcf2wpA7fBLHs
uOPpRRLDQoJnxDxjn05nUNzGAYNIGfE1TWUHVAdLIF1dMntAIyScyVEAt9FXR0el/VMCBJDLYRDf
wypjSB9QN1wLuFXtG5PrYpvCsIHq7Ac9GBRqtWFg95Yp3bWTQhpXlOvIuAHDsO9fzcAFIM7Le9e3
UaJb9gN423JYl0Avlv2+CPfIidr4X/rM28s8H9nQoE49mzn4eZmiKS8IvrF9YIM19Ept3Yv4Ct0L
w/UaImjSGj+p65K/bc4UYMYzUY0jW9i/wDO0dpFnnITpa8xq/7UlXTldSXwj6zwUp/ti/AbC1t1M
9nBMqtM0ciOvEDWfRPnz//fDDGj3xh9TmfsrA8cLahAeFq7X7Rejfyhwu7tsP+DwvEqDEo16GC9O
eMq8V7PAArQeCyGCfwGNwM3BVa3KIY4kiDQNK4+VXCNTLplmSZsNwye9YPLFTUn3y4XghvNLWwsZ
8OSZWgmCDrWCsXRc7pscmWXqW3nG0gkXnxxogg4SnwzsuObcDcrml0YQmKEPS0mrnnibK3UmxbRt
WfgPxERpUh7WyjrJgTbIlbWZ+RMXvRpWdVKe4RjVjg0OusTj/kBpFjlF0TNQx9UuvNaw1ccDsNco
nk3HtTARYvMvGkG40W/WrLfzZRe46cIzXzjwNbz0eYUM5KXivOXg5eDfnReJ5LR9Z96EE/B+M1tR
+vRFr1Es3Nuscd5862/J0PUuN8HAYFKaPBf8fZbYxRIQ5tgtkXZ9eNcCaw/KfTJSA1GCM7s3/AEb
RLIxKkx6POE8yMRmVpo2tyUgXU4daQA+fO7kFVMf5EP4hn38p3pjuYwaYO96k8UGKO9qcI5CFnsb
JKWfjfb10t6Vk8DpXRo74CgbkMjjXw36X6EsYtjOidWMW0DzmfHKZ+hoGPtT8XcV6r7SSF3Yvs43
QfVBtCyRREuYk4Er7UcMgZCLxGlPUQuetKSPluoiQZ9A6DTqMzJKrc45MoQD9IcioqBc+QSviD7D
ZM0eo21CqX67a6FTcfKtoX1f0d03JXM5Vl/XfGdlYEIhrfuFtY02slsrHcHwS3zFb14XADySq1va
qHpSSpmIhv+p7jmB88WkNgdLr0qwCvJOAXldmiWeQ9jihZuiT6Zc3K2Y38X0NfM8vHv5Ax04/Y4l
WGbmWSfD4Fyk8S7I/K9C7OWRfKM0WAJg/c0xHv1/rrIlwwkskRXI2JYwqdolCbB7jQOg50TX7RWh
sF7Y3DyLukfGd8COjoPv2Bov+rCShsSKsLw94+i52/1YUKshq8VfOHSQuU1hW0YbkudOsnZi+e6e
oeGySToymVLifDJBXXScZ7XODGUnge+ikvw5vc9Ap/UArqWPG7OmenFW22ZcMjwyI2fuTsKMMRnc
15ffU/Ae/rTjB7LgZ+LJ7lRJHkSI7E6LKaDOc/5If3x1qWhLK4maJdGptAofKKELfm/jX7Qa0+o2
WbfPbDRHfvpMd3vmXQzwtGHsolYshLKPpFbuq5d6kFzP5Iwcg3am4WhqI1RnFjjKwG88slSVj8RR
27zPSxOhFx1JMcHZU78Rta4abec+uE64PKtlvwOPWK6p3mOPuvyy+5wDFJ/YkplThMwwVmzk31I7
irz75E4XPdde2GHm6mDQGDjk8N4Z9ndhlWkh8RD9uAHTgSNn5dOQaOiRi6AT24x1XCebmZ3jin87
VxPp2Iwq+PJgP5k7OTNmuma7MXDprM4ZPBPG2bCCH9HAxrBmsTcBRL0BG7IkuYK2uMHbQLkT38Q3
lx5WtAleI08YQ9XNresDeQgmB7sjXx0Uo4azHNlKt8YmCNZXaxKFDqLzAh9DF+J+SKj9u4SjYCnu
EPtQwonjp1x+bZggFiAqfpdd4kBoLcjTfBTkD1nU6b2GiHM0RXbMXzPIn8xvWx1+REeOML5GC/4i
7cOwzkMxuXedoAriqJFI0OcGykj9B7Gig4X1+k4NMw8XHs8ipkXfV+C0wI1IRPGfN2hBGk7iVPC0
5+QJX2Pq2j7qdYg5/sb3E7SbX8rsb/+yFLC7HOAyXfbeMX2VO/7kpyuksilitC8C3yhD2ETJ7Eek
vhCFDrZnx5VKDO7L6sZcdeh0qJ3TkkcnwBgpX0x0v5fRxzbBOhrUv4W16n7BB4RVtZAeoxhTbeG4
X3D8Z1+laKnjPAdq8kKaqgdcCObRu39dY26hi+XMBRIImoOnIfIRVn5SKVhUF15ipClVjG8JkUWG
nmj0BftnBm3/e10cuGx/BnpLf+Hn/TX907DHIntQGgfec3xbgPy494G0leuQH8Egb7CD2yyv9LOM
TC/UZyftCviP/r1XiFbX3r2W8RRjQURQ7IRMWzGxtJNEOGgE09h73YdJvtjhjBA8eg9CJgffZItL
103sBvRkYoLEM8HelxQUuF62fE+xnYqwkaO3dEKI5JBXQBUmJOusToF3AV+8vWcOL0zBov7Arvk0
GNhPLnjeGkvhdoTL7hFDJt1WNklLvZ59bes/9wF8Q5S1XL7RNS0SWZKL8ugBS8W1RO/1WRgRoFHJ
soYPJfWek97YYtwbb2GccZNHFXvalWCf2QsUgsAdytPK+WL7pDm+HEnMzLbM6HE61K2mveMV9261
e1zlPTWQnu5qkBJBcr2Wa1TPFEmoZKycPLkCYXBi1UeHSSgPvqKj+SOWyzEaQGRGapA2qH0hpkwP
DIIbMF/1MNhlhDpFdPCIuv0xqR6YIrV47GPC7FiAJ9Bv62I6Dv+FtUrLUjPcGFwAYGJ9HXKbJaQq
c/4Ez4Ii7Lw+i5ZftukiMlh68cxFz9rXJDRKmk5qFD/xXrDDJMCaraMCPpoCodaaqAZP3eM75mAo
0D6kvyA4BwN5bNJZdi4dmCl65tOPsMDRN9IT9mmCyRx1KPtgi1zTpsovTN1UueRj8Z6/AIfQrpeN
sKhBuNTIWNtXKvGJuuu4kU9TByCY52gLcuipGs7XlxOIGbHksoOwH1tngq+qUkLWZCOmjDytGLDF
cEtwDQ7bd3VRbWiRQOylIHnRXvuesnb1GDxIBTg+/iLF+1GjVANMoLR39xP6pIB0P9+mN7pT33oB
nwik6S+aO7vVuu2bO48GhYeyOoWYZ5oFJ0+tIe3/UEL5XvX8nAYZxKanC30/FtiUiemp75D2fM7D
KpMb/Lnbfg7FH7UVvDpjffBkP32QApy5ab16rJsOa5s56yZhUqfbamav+rf6NA+CamCotRjiIuFE
pbk2Jf+BuwSdXTqiJ+cxnAs61kgJdVnrzDYx2AzzXabIXzvNN9IPBnbNgq8snAE4C3fwj3DOFffH
6IT99+6U3tHxQuAv7qSPFR61vErE7ugyO1LFLXr0sNvcW3PtL7HaURBbYJDC5hISvu7TJjKyL+S6
oIBXEHm0kwtTvgr5NadZYPyxq+1+Tk7XyaKXpdBFYtxs20ZdOf+YXVCfy5kLnlDM4zs6UmmtuIka
e6njgsOVbfCwO1hpcVbMl3ZX9+iTWuRfhRjdnKxqzBx3d3uX7vEcYeJdrk3mBFjTc3IEGqSBE/Rw
Dav7aWkyzPhuAbDMC259RbhUVcazhaRULUyvVSsc/2ErBntIkNjdDw0EOZaiIDkqUn3vXt1Ff9tm
rQAUJo8G5sPMzIN/d85zYPDLzk+/bBn315+j0ezOQ7Cl7zs913MfMOHlIx8wknoVgHWExBXp8KDi
bhsVaEy1T0Ot9/mYvge3256tvQym0zSupJ5wYeWz09P/ouNOBDzBFZLdn3D3jB5Jl/3wszhSJTs3
lyu9fFYAONCD4AGzKUprCAkSbOuOG5Qs5CNL2e1jg4sZ/gbi2228+ZWqkZR8g1lQ4Q3UHgjWRnaM
HpljiHXZ72cHDT6Ox1Stl1QszLerhF6wfXCf7BsMD1Or2/ywH/NEHPGtiVxZI47cegdZztL4cwKI
4FqibBF9JGGC+OIJresptdVLP+hC8CGYP+WOb5Ut9gOlQjBfeaztHqz25V0lFJVfOiKhKYHAvhFV
c0mEsfXE5mxmjJU9/iI9DckfaNhuDXo0Qa4Yjy9ZdsEAuSBg+5ceaLbuN8SOGBMEEHX888dsGjFM
WcUWAZHs4wYoY1YoGGe2Id0qrcsGUBhIO+uaYp4eogouGgbAA9H3nt7GFEd55gEPtPr71f4bH0lT
M9ddblUAFhb5TSjpBA8cnc3wi/DIAdQHXR3nA4FbIwQn+eUTdkvotiPR8l8LQFQmhYYrUsURZLYi
VdGC8yarnLw4dosOW4ivw7CT8CYOC7ddmRTE3o2k5BiHu02U/0iaXQtJJARCfsrkojx5aJG9qZni
O7fliTFx55sLN1dNOzSvJK5ZpfQ4jt6mclcpAntdFpQomBhGL2/PjHur+vAU3/2Q4RV+6O6IGmkb
ygFz+iD2IyPUoeidzZW7FdEx6Eo0wfRCx5Z1PHdt65ktnYEi44X1QKdXwDLbTjpLRukkZDyOZXOe
N4Hh2l6eL0TvVeUwYuLzTJ+o8Z7nVSHlhlDZeEKOzAvsk8nZuxjrhXgPK1Hvogd87wxyRZ5yT/5V
flWPg4mdtRreQ71Us9F61NuZclUITRG3Rtp7uE3YYtZjUUWg/fJWlPq7pu5lJBagWACg5Ow0hg6E
FDtEZ+zAu15Mx1NiOh3Fgpz2wh7GYhIFK9TEbJKciA8niw5K+wVGXJEc8k18ATEikJdOO76WjqBt
fWmzEYL4CwzP55GyzK94bFStQF8qmc72JlMatWd7FZlFPH83banVMrN3atMZr00poP6wnXf96Odf
zrmeOPfGcLd9ntufG6r3FYuSPxR+G3jujXKczsxC1WJbeoAN1SwOy8M8uJtlqXjrfzrO5KZehn4r
ZwZUnw1HGTHRRuixxOozmvql82Z7s8JUxWnXR9AlGLGVz5YAZ6YGf3iH//eiU95d8LKVoJGAwjJ4
zlx5FxsJ2GVoBOfL9ToL8s0ocZb5vKXj4n/+yc1G62DudcMrEDRLCPF8yOzNZg1GtpU3v8MdV7ht
xEOYg0mkQm199EBdQowLwhzaaY0zWsqe11NLGCKkNi7kZxEmyH3uUg/oMDE3hw/u93Jfk5fBbp+B
AANLEwMMTJ2qGqPdmcjQbxw7DPtUu3unHQXnBXfcRJo+iN08BD1eiZiXNeNuUaoLFHieNzJpCJUG
CnK2bWGXGA2Zuv3SkTFpDOR+YXGpPT277XreRKsIwJEbFiPSh9cIvyIlksj9i048/W91FtZGsJqO
0RnydckQw4rH6Ge9XilsjPzR/DFwUvEkVNx7LB7Z8Uhmx6QTNbm93KzHUtmfOzC/c+7gNgWMSH+3
1USGVDsNoxBE/eWTxKGaWiP5SC78EqMXBbp0Qr2ddht9YH1KR/F5q1gkGu56KjyMgihLv4o58MPY
NPWq4w5n7Na2ytT12/NexS/NhGGe+RWMtN5teD/i8rY6JDZOBYuegvQXiwfDG2CdLQgdnal5Y/tQ
TM0nU1gFSlxhZ2GFE6HeD0LoQj/cCL2vhSfmdJSsT8A3VZn13z/b/8KIfLQTbgD/9Zq3yLRCPcRP
BNy1kftuR6WM7oR7guZCOrDdtmKXJcb2HelikecphWgxm4CbPFiUFohCQPEnHkEZImpLdP/IH+Bj
E8Nb+ydn//RStN3NmR8a35Ohsgk46UNrKAeQWHOEiUc7tuvQjVTNqtUWY//W3Q8oLQP5d5Bh0CJa
xN1MUsQ5c0O1Kj+H+/eVIAlSSZMqQTcZnODUaj8I+CldiXybclpUw9XwkGsvkCRGVhIhYu5ucixp
dTkyatfSgQyt6JcO6j9gG8+y2F3Zio0xrenC5Kqkplb1ciUDMnSWdYvEN+j0ZpdIVQNfZhCfMY4Z
wH2/cZZswUleAWxKSLG9f0oJbG6Ke/GO9Y5L81kjIQNJsVCRaXLlGBj7csw7Wbo2KlAIB5u6ZnDB
DMa3LKqYQgk43+jAIaNaKbvT6bjMIbi7h5XmVdqhYJkkixs5Cv9XSE4MZIXU1vf3u56fi9zmUIPb
tDg0rBMC8CIA66HSmRlJV0b7KmgA1aiETfiRtDg9GPPPxweDBExs80NPKUS8RCX1+yCkSbOs8lG+
fn+D7ltAyL2t3UifnbFMAQN5alj4vYpi9huclnaBaFzNjve4ZRY/NM4JfB5gHh+r3zk4vNaaSwti
+2kQcgZZn4sNVuO4d1GBDl7JylIu+jVdMPoH0KVI3Uz6K1IojZ61gJ2ogTOgRdzsX9t3yh2TguW6
k/6SE2dQPyNxHZoRnfx4KQlMVTkBMTJLxWH39K7A3d0naPNZxv7WQ7XFSYnHlctO/WJnvWjHuKGV
0PuBytz2g7YS8GQmLSr5gSMPeTMuAJwdN4hjCXJF/+rNfzPR+0oKH3D/ieyPaBZlWBcSE8yzNiHZ
vLVBXhzgvPdL8Hz1XnePixFYibPEAKadfq9s5FTBDbJqVbuLUsRGiBX9rEvRylRPYpQkoew66c+T
n9p6qyqlQFXcE+oHWQJu/FoubLU3FzlkP03d7UOovmWH+w4Q2rY90/SisHoSjgSi2mLQSbviMAjH
+EGVWPgmtVARJEShdpDyFLVS1m0Ba05SOGEZoZtYGIMI2/PE/J/C64U0Hcg0dRAg3ZvgQqWo2r0Z
hDkAIaf3LNBlgu2n1XGnct2DswZOoVYuVyScBE05tzb32RokTHeWCCc84fapMg+4DiuGKqZojC/5
xyFinwEKps/u1AFbbIzVOpahHn9prnR3+x0oNbwuW6Y2hTBj3bNmXkyOZAAihRBa9jcgAfQbx9T9
NumYRWT8wnzmF4cRrnMVti9OaMjclclNSuMCOZQBdeXC399PQN9OuX7LOpoxlUCZ9O2S801bn094
Ymf7Q8VqJqFVrCnQ9EZVk7l4t9psJvxUMYrqCRgeYVxSdQkm5C8q1XBKz6MxkcTP8p2Km1H/1tXN
+tOSF3PFA0tWi3iYHGn45xRBeZgVfkVTneJwtLAnv2CnRKNqoRcL3GYEAFamUCe9tqJ8JpHyZImI
VtLYEYRx8qLzih8DicPdsmElZu7ZurOTit67DcOPN364ay37zgM/iZeT2wcdniFeINlC1oS5ZfjR
h8eCIxct5188X33gjPBEuOkL/2mRsFgN+rfGY88oKAWD2aaolYgfzEPBLb1KjmkQhopTY4TRxWO6
c61DueI0fE80cvd/IIO3osOK/qOFb1u1vJ9dTplR+ESliz2fxvpOREJeZFDCl5MBaTjfv23sZOiB
bB3cmapOP7txVjqDOJeWLi9tJXkGONTHfJWP4aZ6QO2u4p1Gi9cRWyR+wvK0nmDSCpH3xi8dzqHS
sbyUwRlgn0DA6T9PnDtTQEPOWc79iqAKDAuuXDd7OcGhaSNjpKEG2J052jqH89hvW9F9+n8CM17M
dL3wVJvamIJTE2/HhVBp0n1oVgi14RjVXj8nyd7zq963QFfGSk/DSSVx+cf/yA7scwBuwTEL45m+
V+EgsmA24HtcI7kp39iTBXjWH0/WVxHglgYayD0X9KjcoDEUs8Td1Uy+aQpbS0XVMcJONVaf41OI
ox9HcgxsQNlCucOI4GgMNmd3YBQy2thz0oE0TgG+z/0B4p/1C4ohkwuT1z4jxIHwSQz0GMiFsanI
G4qEyJMJ2vJ1Qpq170V7M/Und1gz3guvJN/kxPl/YHS48gy5ddw/qJvw1qBWPwdG3Adjloo7oY5d
4NNlaCQe6Un0pkjqP6mQY6M0M7vbBq4D/mbDlLFdSQ/3yijFEn3A6tM6S+Fh7whSmQNBiRQ0dHFP
4j9f/9B0ggczYJ15ZEiDMy1JYcaqwV4n1Xq7WIkyyDBcxJzF+UmBXskjD/ivrLfe34wRXruDngv3
rwVSQtaoo2hr6IAqMcOZpLHmLICbn4EQ936v3xxE1akbcIv5b+DMWSohy7qX6wj9py1jUNwXcquH
NPlvUoiFPfhWIMv2f5bkY+XbRBVLd7MSWZTFRzdSF4M3nPaoIDst4BDIL6EfGkddlZHjdkZtSUaU
zuHA6jjTiH/4eEtQFX0Qe43qpVGfrvQ5lLaPQpKP1gIub/cj6zAdaywmpWiObwm9BLRbGOjXCUX2
kTKEPXvaHeaZEakkfDSRqcdzOArweeRx7OCs4JgG6qr8Nb10mIVxzZ9nejW9AKNci9MdweuddDuC
481e73VVmKjFd0meq3l5b/T+diK36wp92CUtvYkVSz7vYi+vihtguB0566nJ/JfJK8TSI6k4/pt6
1oLZE2t+dznvBM1cRSDEE3r6QK05sKdyqOCLBciW7grkhY4eGDZ+TvvoXkCOzPfIqcl7JvEvG32h
QALtQ0zREpH182ccDl1WHmuPrjIv0LKnnVaObH5/B6/RZys0s2WbLunyaH2GYWBk2Zs+cFszL6Fa
ZDBCJBxC25ncS5VAxxuUPknpcsCIPOH45Sm+nQhDAB1kDP2/G8fiteu5wqPtRScM2og33hJRvRLN
cPmY8GceQPOuBVPn15Ur8lAW+tq5syITIm6at3N997Ew+yCBKtgiZalz+chBqUV8w4KcfSELIXAB
3iuUtmi3/GkoWKIk6V/JeoAkR0tiUuzeF2zoYT+q3JyeNMOi8muT+2ivqEtMnFmaouq++QnGS40Q
18ZEaXvgcOLAiSiwA9mxmcL9qruIFE91ROG4rodcHBgxlqIbP5Aoaw2FSkF/ywHwyvw+gi2C1UPy
W2uwnBV7aZJjckAEyZFwvnEUNZVq2RRUrujIzuON5UvOHEUI4r8uaYS8uQBDS7pT7hvLR0A1BwFZ
I4NmEdz+AOQBQdK7yUO/f1JrbhKcpukZPJuyDd02cE9tHE34B2eXMrraHkPOV/rop9ClhSU7QDGz
xmUVi5w0l+YsHXRbtUtag/OE9JpbkX4zhpBdj8lpOSjZbv+lGcbd/yKsw8TytQDdpyyBgM4eRUlN
eV3k8gCla/myOYb5f82UXEEP5esmK25xR1DEVs7tRPEMQNAVBDfkf6P5WruykUuN2pcsLMoMbqAa
DfTtU/1QF8EguS/eE63imAPtg00t1s0WGp4U9+OJs+Ui40G3eN4cqu1oH+f0+h1I05lq87hS4vgS
AonIAodQFYf11bKgvDiBl9JFvusTgz3NCcTMNH+ckzEmepAjtc/wkfQisxkC5hKJCMvv7wv1jgHV
ZNOBhWudLfauFuIEpyVY2IFa4c/WhS3fVxYywI6XMvuxtzGuLnhVSU0vsoc8RlLLJciPbXkNKGlw
PzqEzQfe3n0DioW3rws+HSA6Rymw2YlnumaBO4kDNivXGBG+b5v5uphEojjmRRP31C1yTRH/rx09
9XxIZEKCTgL0ADXkIwpN1BG14iJiso1AF63aYuhZiFeVEa5JHTU4V91NmIODMHKQ8Ffv0o1YQ0AB
2RIkzniDIPu8m3suMVpiEzPOl5eIR/DJ4NS71lQQQaSkmTzlHpN+Px3yIEVrVdSHhrFDpcXrSRwt
ElIONa9sqbYjbgsV+XMKMBQtWjOXi/fOel+c0uFGBF8ibDuDFfIiS/pdJiDpEwaY4pMLC8jGUz7q
ofZrovRiRhY/mB1g9Q/UGjDj6u7F11Z3A7/iksiTocXbeuhQj2GhQu9PGuBh1fCi0z4K1M7W+Dw3
XbQMDynr9hS+9VNtplrHv+vFPkPI1yi9N8kQ6rPnwY08Xg9Vh5dCDEdB/GwVGtxxnbyTpjXLlcoT
Nfnye7gk6okbRvi5xLWplrAvnk6b5g+ZabZDaLpitSsIoXC0oREPY3413yt/pIG/u1lrUh/lpqsr
V/dzVtqs08vGrkQ7ZkXsrjU87KTxscyMlkx9hf0TpW6Xvmk3Gffmvi+frmF7S4HPmqr0M1R9yw/p
YlPU8leOtZfYtxXsjq2yJRo4sLi9A0gPWfP+L/VJiRUubcsp18KuI08hJdlhgJeiavSLtxnnpGC9
OZzK1yOPqi08ABB6KKLi0Rdite0rNaZLEe6Dg0ZavtN6qJr8lydUiuR7F6CdHbEoXtt61oXyoAR2
dyx+FgzeThcJvTSWakXTJBAOTuyDr06LaPk1IPHFCF8tv+8eanvvWaQoa0flu9xdRNtRpxN715vd
ykAih2JiT63kjdYkDXUdpYzm7lGHZLey1U5qiBYRqfkyEILkNWPupSijRgyp7e1Zx2oT3/5676Ll
QN5SVZLnLVRfGlzyCkgv8aAO1cmzE8nMjPdoQx63En/SZBVayZdXDaW3DiinP2HpRrKc3yCwqdvW
zuHyEaJGkF73Qe7XAuy7z9FCdXgmkOjmXWBPfe//7ZyLUo5DxV3EnAuyLPQviczD24xo+cY5lkhm
7IGEfdSdUA149bFpoAwcJr7GLmk4yL3K3FDmxrQSZuR6r9XonXn/HCbls+HqIMAO/OM5Drq0jue/
/Z5DIrHnWGHksJgFNkVacGsbb9Kts+QcmNhp2h6pwLGLcw2ayICnQg8JZP6miB+7kGXnjwxWtRh1
ijc4bq9ZJB1usLZ52pGvw+8iEzzc8pDKMBSIFGokEpKW1RmHlkR42GTkFtCQmwHvsSv0zOIvAL4R
H18pHtTIEMxt6hf7ht9/QIdj9uU50cQ6Kpa2uQ5iT5C7CxUrwmhEqvw6l5nAtZ3DrmHr2AEqAVPF
OXgrP71dHwD0CtW8a62R/07wHEqExc4ao5nrDT32+yX/Uv3vMzfVnT9USHTdjtrEN194LgD8v/T+
KIjty7qWajDOgjerfOGWHZm0sTjJlCLilYrcbLvAAoD/hQ0Nne9utEHESEcXn8B7t58vMxgxe2td
d6PhpJQGN6qkt9SiDZx5weP3uU7uUBcExcHlOFfi+JJr8gHYazF6pW6jaoGULafY9Uut9N7nhiSA
uUtnqBrZUFT1xakuHidfrQUTbGQH6oOc//NwXO5sJsBkes3vnptFScQat5z2vJerL5wIwkh1HUDm
92qxnsukH9Mipdx8TXC0aU25yhkTaULN17cHmBgJrfNvb9EiWSmpcXabzqTTNu8hLoctgybqFY8P
FgYPm+GCuHvvwlzy8kLohp7oSoM6M51dihwBqfenXx0OPUkj4ElaLD4UzmyEPCepjXf2W0ST+Mnl
lauqt+VBAitMQi+pB8Jo/0meKc0oBY9i5MIseUS0MkjKgC5zxc4bKovcdNIyjH9ygugVA9UcD8zs
bzb2u/r75Lj79WYdZVHixcTj/Ucy0ocEfFvZnhHDfthF5GdOzW3El6pOO3x43qCYueay9o/degPz
f7W7KnMnBZGNTGXQbl6O4sTursCCF0GzznPdo4msxvY8omfSzaypx4KbN105aogcSGCwloh+0puI
/iEP+z8tRMTI3Q/sJVT4YHodit0RlaYJbgaYDpDw4qwcqXTKTJYD/qqsF2KStHsr/lg9lMmHn3iL
KlRKPl/F3EZkV7jp+zRe2iqz0uo2hhiUcR7BQleE0aIiqWYCLLo6mPiM0qbxjE3zRa4S1VY2Q0JU
Cne2JQ8I0v9XaHFU6I1o4lyVPCqjmNcm48SMMc9d/dcQYc+DsLMmz7xmaZt58maO3DgKchRygjXI
9M5f7EnfSqWeTlyPSXzViOtDxitvGlPZf+5WlW4TcPrhD36C/cwifiu5OtywrgLLeP5oYWvtTPfm
k0gvkP2x3M42L15cKTfrQEvTjiaZ6NyIx8hhQLJ+wcoVUxDJEscTFT9Gemldhxab/RjHPSb4iy5+
CVrSciG+A7q184C6oCzAyl6E1G4W584zgIyEiAHW5OfZVL25OJxDvO24UN1ioPFBXPloHaG0rjVE
9FZ24NIf0wUqaS78U1hmUZN2QE8Ypy00xoAHz8GhQ7MT3PVBg6dqWqbvUkk60I5ZnoyjzlGfYpYM
sgXbdeHMgidoTYrVoGxKavSLzoFUSnXPbcPpdq6sG67zTjYMLwujhoXzpHez1ICeRS9vZP/ZRHaj
9P31Q7cVIhDRjcTfY1jAiK5r3joAWBjABRV5J9O8ogYx3u/oCH8/DSEoF18m4UZ+h7qBXzAL4puT
zar4BELcDnM2rszpefnob+8U+Ew0gK3DPZggCg6f9ZIkfNn967vBKDRKIkEo6BSgEyJkwzOGwB2o
NEFputF/P/QhL29v7HZ6TErQALLU9Yvw/eug8FCDPGVsPgR54PyIAR2FW2KXqE7CDLSvO794Utff
L1HbPKUZaeF37DO4ThtyVij9OPf9If9X/SOUbBafpzu1coKfq7ynZ++iuzoCV3uPxRmDHfdTkohk
PmmawL8Di/rDqv0SHKotYmi4bAK174j+JFWIIGrJ2YgUMOh4vh9SFfm1U45uyFzDAZulfgaO+9O3
u3Fckqz4hgRhsUthHd26OxmmDgVn3xK7L/z6EHBkTljqKsMxGQzmYYU4c9cenVkiC9QFt4RDvOcj
vT4w7nu3bbc0nSX/bSefCq/EqIXEW6NO8g5fRDcdyHO/xyY+sAEalSrlPVAVBfuh/wOlEJUxrAoA
lACTmL7UqH8djzz7ImIESOb9AYUKiQlZ+k/ubTAGkVq3YNEZdM2zNxhczRsLDoyY1qfDuI2O68Bn
lPsqWc65oTodxB6Oyi1oq3Rf/LLkiYRLoJ+IRKjoFJwXuKbkvbM6WUBsefYLOATus3L8ZLAU6Jiv
cmcKqL1skGPu7STYqrnoJAy/tyC4L83O9HiuUcf4ExKrHDfJvO8Bf/dd+2t5ldMnGlNTwWdLkHmZ
Wwtw3SY3wT8BftNWJTlQ3LxpZ3/q1b7SIVdhVUQdOJ6P7QAU+JWL6zrII+jRr4jVeEIkjEk680hP
udCv/O9rz5jfdOwNKgPEj65d7eennIIqcCC2go3DrFK7eirqye7fTVsyQm18TiXLmanoDJpFwopK
jY7Z6L+hDYVZRx4vVZBeivP5uGpAT4R+v6ZVV0U9lx/0Sn1d4SU3jgvrzo4CZf72WKlkyHcv8WrI
DM7uih8cmIzZSJIf0bdLd1LtKsdw7IvQbGmGa50XUOVLV2rZ9FVk86cNxxG1qoSJxyBqzF5PLgJi
dQkCApB8qy5mGPIPjyV+WeZU1xLV6maWVip5vlEXXE9pF4RpLk3GjFrMsNse1qAWQH5mp2qaQIn8
38ue/nd3YAqQqEa0komP/+7fpqJH8JF/+jvYmAuPNjqH0mXO6mm7KQ8vOomD5fEyXoDqPOcg9ZEb
ANlqndWwd8qGKFkLf2IAjY1Ci4sjhE/nOl8rz9wxR2AmK4J3rO/69f+m5nANeME0RkjvQzkNkrvE
d2Qy/H/bAs9AAybtJGt4YfOUt8okmcNXGzVD5/BxXvBYcgQEQ3vQu6bKsttggGMHvGghpdir8CDr
yE58gwSH75PD6LRRjuvG85S2XjB01BBSs7QzLCURyFG+aSrIbih+/pdN9RxpI1X6Ag/psOVko6Vb
+x/FU8VgA9GsAH94KK0p4gliUAyXxqxvAXi1yg+Dq9TNlDCniLEX/MFdBZwvQ1vI752p9tGXGnWY
6QqVVyvy6bNrfKZBeHz4iiGfs6HzW7oqQTlxm4eeuRdUqEdNtWJsAfw/l72F971D8pg+yFydOC6Z
PNO+1w9Ow8lSex78Q9nmhZDdOykjiby7ubarfxCG4M2HWF/ZPeFBQKU/zbdseR+2EBI+dJvY1jQI
SPlV2uIrHascwryBJhELkYwOPG3uWo4Pu//PTTc6T7S49QGeP3QnvPlH6jQ6TtJJuiupQ0DWM2Le
dFcYtI4Jf9JL8InC938FKCDd4OI9YlAw1jksbdbRhbk+a61pcEEsxE0gXusUqRDCfnsghKrMCSp6
XHZCYlFMBO9qc/VkE9u3c6lVhB5Cx1h/DZHBnwdFdNqrbAFf8RLFGZd9GVK60hCY+ZPxL36VvW1i
L/c/uKzAWxaR+T+sh7H3MAISHLDH38nSPPgOubGuSGwu66DDpVl8l/SyLMKPp/phcCnwZACEUM6M
+15O2/YYxB0xJHG6hxEcCI9GcNvPE9OFMt1VokMsLsBCME303IRrz3gSnC57nXEDyPTljrHkIMuu
ODtSAhEBWVCHPyzL755Xz3rM8/zXHaYVrvrzqOXhFEmei4No5wsUZa2aDxTOcdEVrB6YQ/TtWAbD
XMCxdfnfn8x5P5bhny21EyUNcNStGYoGSvmE+UGnwW7n0cabLYHBSiqurksQL3Yp8KrEOZpHzfF3
cgkDQbxRtcM9e0DeLMiwkyZuGZDx2sezTcr4a5VuslGPZYE5t1MtF4UZufNRpouOJeDeEoPBZVzo
kBzUK8MvAtlkYXeAMsmn1MKwCML2rUDiXkUqfGS3QdE/qrsL7EVjndzckBkwEYuIuMSV3v0Wqr0v
RMl0CxCY+LTiBM0ICxc5iDtwaIsF6U1l8reDmLAoaPEoIOb4FDuQIskZV8p1WY4scDoK2I13fIe9
N/wh0KhRMWMvtgPSU1mY1lq+7zM/ydD3bge6EmpPuRlPKbZOfv+aCAf4P8Rmlzx1+DF1KdHBKbV6
9/EZVBpSlVLF2l3QdoDwNTsbTzKWG0lfbIkXngj5GLVq3+s3PsQilbagYw7tg0eP5dU1dEXzADFm
hblTP+mJTq47fGoL+VzAN39a3svgF7Sj8B9GArrgMUdoMA6IYjOCIXdTQmkG+L73OM3vYGv79AkM
wVGDhDC+wcCgtT8jGc789l0LKhbP2nczkXAwmIiVTb+4GEQVerbZDKzR3Hz4r/f/b+qx5rS14r/B
rUsOuH0XKiYNDKxWbN9XWqOeQfmhWlKItZ/FT0CaBRdJ1HHDJdKsoEL7/RIwVgq6lEjAj2RTKmkY
0urEgjY44UTjQrVipTIJXV6yalS7m05pNEelNH8/vwYuxdpmjZYjP7YBe3DB9kLe3XDaKzwuKMCU
DttBrGCKBDf7V7UmywwKzALgi3ifObiDW2AcJ3NdM3iRpnKSPfEXmyJVSNi0bATnUKpEBfPpvs0S
JEWPhzDCzW6ra13x0bdshe788mCqv9/5PSoddLaPViMyvO+MyK7iqzkRMkgZGL9fWMmYfAxpd1Sx
Qu6GG0K8wFUSwDPX52UrrqjCuf5upXiw6OMtZ7g2WYhDAPJTkqqqiINbhDRGhL15RXiDQJ5y/KKX
tueFfp36kpABl4SpODpjvPjkHNNQqP9f4K/o9ZvafAdbhp5qFcf/gm1dL4HSFYW1OhUJBoXdHDAv
Ze3T7A1OSsNZ6wFy0MhrigodTADWuGlfkuoTq5pZBRscBPmUWGw+sYD4I/Fa8T6UsuIlVK6hYlKI
rKWpJkfyUBOPbNiuGNOj2JjDD1U+Xi+xPAzlfnyNtsvmBm7alwH8w/iZryDtOqZh5y7sja0P25f3
tQzAaRV6maAqcZXjnfkxIWv4GWY04zV+1i79fiYr/dEUT4SHHFXBy7l8twXgtxAfI25RGafADxEL
L2f9xemLPG8t99A4P47ON6eudrN3t/gMJrPZKa3MkxfyjLgUd6WWz5rBamvz/QDMkEl6gSapv43p
s6r5mh18FeNs3GaqnU+Roev9Jzoj3nBFCfWqXct886kzzAbGjLedwPwyQTqLg8KTZblFussE1hSG
Ryb+XBwYMYxVimzGfor5pYfx71X4edJRc39466F6CfA/st/gaSzSgPSurATb64CZtt/biwpPfQ3S
tPwy7l7rJUegibfCQosVz/CqjP7ejWLPYkJjut5gMXNYsoKtt8gl5OA9eYThzL/ho6JSJIUgRExr
k5Xq/wSvMeuY3eLAPAarSwTcR065NBENmVVhL1DNBl+zs2Tr8B/p/S3H1k06v35NZQbKm0P0tisD
5u+cBoNygHsZ1UoipRN4U8jL4Lla8VvYdz7bgkCAyZMtzMPHaV1zMDzMH4ocN920Roq8nmW2jLwh
LrNrFzEwj4jfddQQxqLe9dpJ+bNENL3n/7vKDlpdYTj0tQJw0qegzfsTau3mtwU27sfaiYS77sg6
gHFdWUYiCcJ8Lqg65lDr6njoFmaR9aHsodhNGXiQTUpPdWCej6A0GuzjW/SsNKIJHy99qEzlYenV
TcE+wxNq1aUm7acYwY0MHl4P08UP3YPhlbCVWcYezMofwAeYkeu9zHZtukUddOt2BSrQN3KRAFK1
Dtg0WiNSa9BT7BaT68Msg32KLhGAb0Wdssvfe4ZyWTDqusb0qIy71vlt2QKdFJqBsVsoLs41ARwr
s1G9tO1UUB11BXaRWih5qqvMzs9Gf9p+pnsLCEGSdOTUxWSjWz4TdzjVmCAxCNMI7PFsLrvyMT99
eHF5oc627ZQ70NZ3qzwPYUacmTfvv9nF+fGlrhZxqVoG5v1NJHAsuibhrWtwv/4jFrzY4vWevvXw
QH0WaSlOTbtlFkplD3d+n/lKLKMsMTLp686IcTcObdzItLe3J8ewE32NtT+9Q+5gb9YuPVw+0EXG
IzN5nZHOw1oHxOh/75hYYf8XsSJEOEm2Oqnaedn+tlCFfDNQMZOdRZSTjI4SgFziI/ohpMNLqIBi
go+MN9St8aOdc34v2aozuvqWKaQug/2bU3FUqnGF+Mg32JZv3gF02hIEWxrUTzOns+XDUVKjLRcT
9i7IZukeC+64khFN/9HLGd50rcQTtv6o60lOa4CxJKv0JazX7VVOoVlGe37UIJCF71khCGyfm4at
s8nODxKtf2IJfR3Xgul00SpylhdEYwCtDBpnVRQkxRj4v/hRwy1NDsdgWf7KpwXtZ5zIv3A7miRq
ES6aH259C7oJcmv6I4S1FToscQWDCJIJkwe/BFLy40K0zF6gnC6ZC58neBIUohsDbHwjlVtxMydD
sp9ehE7AbS/f2Epu9tDHlS356/GitP19DdHyMJ5cgUzq0Cc9cOtzT0rsFMV+0ji0RfYKSrp54Wzi
izhuCIN0ybzJtUIKxWzZtCkVVznsQSwcTlCYT0cbh1Ah+8jcOTsjEWdBqDI7NqcC7V1Nm8DP9t+X
DWiYTrpLYu5AFVdJdjzASO8hGfYrEGSxnyAwU87KG3ZJ3BKMPVRKq+2jV3NKuCNHYi/uHzCLmLsC
qXVZfXSckjm3oVsplP4MqCN7CXUMQ+FZZ/0T0ONI2mKAxdk/IhJSlO3E8zEZaRwY49ulUYY6UYcf
1Lwpn5QdSixAAM2meLSCqCxPbuf7FiM6fKYTm4XlztPbL6q2qUxPyO1hPOhGTdliOsuNKgH6i2th
XfKrrc5tZD0gcy5blhL+pHacL3qDLWh472QEkyUEDPWGxAm5xJXLfF56aRsyeeuVjJynokIioID8
2/CFuANsyRN3dVo7+tUBv37icb5TMJcr+3OipL4iCaEX8c+DY0TfV551kmE95zR+TcZFxIiAEeYU
yGN3cV9s1VXqWr7Kf6gpYnW3wGfGq/2lko3JHgqlbiYUrXT9nTd3zjaE6NO6wrHxZLiIhSWjobh/
sAA3ilp0qJvHa1bEkqHYaYuHoRMwSNmLRK5SfQIUBNAa2cjhC3p44AEJk7x5lmRqruP9F+sNVOko
h+PcrmRlfEtr7xgdPEuiWctbqFAI98ZNzpoRBoVwijoVlWKEC055g+ZstGbGZahY88awurgAs+xk
tt8uWB+r1dndwzBHOVuP/7YJWqnsC5RNzqHY/Rh3fDJnoB/4RKOj6khwaRxy5kxBNc/JhWkYT/TI
wSgh2kAZKmH1Oy12kSwRXDsi4cidUSXn1xgWsb0m5NNrBu8D8mCUFpEbNrZPuDegCi6kW5NBRNB6
1/KKkYa5d46KCXHN36t8qmh+VjC6+yiReJfEvtFiiJERZElmdIX0oLn5Pmd2gnfsz1GvghpyYxSK
n/hBpxtlAouephMVVIcXXJSXqVEcUsZqdUOutZIGyTw2tCEABmrg+eeJu53BjN/PHXuSwhHxe3/Y
x9sleak6HKqSbx2hEDRAYZavkgwxizBNzizA4/NTde4ofiK/5wyiUzndBMv9l460djWG/jwMHKcq
dQfUO1uyLYUn9/R3UbXOJy6tBUMutPmsP1j6k7g6sHxecDNFsSgopNep57UDlEz8u/2FLaZUfB4X
xELV5jLDZX203yqYwPw8BCY64T5FnOBRtntYm5voNpCX85JYj/8poxoqSu7m4ygWcD6OEhfnKNoI
eF69Va74xkcyJg+nbnLBWL5LjuQt66Wn8qThmZoKR33JN7yUuuzxYPAtNsB8YbvqLf4Lgq9fOY34
8KMknOjRBzpBMo3/F+/cZn1X7q1Ec1Ep4qfWoJ8Jimqk8HjHTv60NQ9IkNZKqLiu9IP0Qt3ywgGz
VI3iaa4JM4RoDRhP1Vl7ALzapYDqo1F5w+LExYV4IjAONvmNmt8i6AIlXmQus0cITbZlt+Wyym9C
lounqOnn361ZnfRPrpR3QvXy8TFpb+vL4yxUlsvZvEPK/qK45rNHZfcS3Q9RwtYjXZd0QhKrkUQ9
9JLCLRN9qs2LV3RsRYrMv9dKl5AqzAH5Hi+fYtEMF/kt44a8xO4QbJpBbbeBe/fxXqUCKPtxaMbg
4kMgIYCdQ78SzmRwwLSuJpkBuMlBor50fA9xGl7uup0dzK6qH4Oz4vUg+bbCv/gA9BrcnVtTbjiW
fm/TjE+RXp4ME2jdQ56ZXkjTXQtU4rM6StC27DcHfXj0uR+4stxt0oZ5kWVuIkuIPZsIJqcuT9dS
x9oDtfjIIVcnQu3N+hXpxvpxxVeKsgujskjqIO9w6jWUJpswjl0AM0qBSKkgUd2E0i140PyaSOeR
GPKOvN02O5zQ/Sk7TMJMpKRqd+kFI6gI0iPIbiKEdLb58sQDQZafnyqmKnEAuCvb7KyrAPdKiAb2
Y7yD30LVx8KZHr+x0FeIdhxplrj+gWuSKAuehrx9O7/+dlsUbQoy+rWt8srBFYJb+WHhnn9Cxs3L
3x0QQQYZzfRUdbUMjZJ3va6cDJ7ASxzalc752EaquFz1dZJJ1JxY+6yI5CjFibHLpnf2jponZZlJ
HEXw4uGfgIn4LCATJ0yD/shOynrcEP5/0evSQQ8eTmSbwNa+hOTtXZxrHVfKdmj5RJ96Zn94H/Io
6zvpKxCxeFP/sJHgpq57OukceGAEHi3yEp9UiTb3wtifE/iGRUaSd3m/VQdMjuwJC6kZ9W2zNQaz
zSgIS1hCkbza07EApn4wlM/ZTwFwO5bxpW3enNfpr4v8Ea/AS+0nYtMrKHLDqtJ8XzmIOlxPMrfs
25gBuA7MASeAVCOeyyACGw2A2qLv78Jn/cPxdF+GICa99nTYmt2vnCPBhesMborttXcoS3vrH1D9
I59pJnAPVxvFgLgXs6mmnxp9mdqpNquewHJluoFdk09uw9UHXiisQDI95ZrrV7j+bD5mGiTpYqjY
vDqcqJWwiLwDCRputUNnltnKwrgn+IenSZNl23LCuv6fn1Vi3roH2z0GSvlWAPLQVL6dKpvLNRh4
Q4yJx/FYGByXPNSs15mrSHGRB9W+hRcRnliqDtZMlHNpuZ1yIsGJ/mQkyvm2DSUoBEYCNzn+pcgh
jkZ8cirIn5zUBXwpl75UPSwSYvBlzvsmWYi48SbaDIvxhxbcE3tr8y4f8nY/JQnYNZGPAnyFRYdp
psbbydsUraU1cI3Njm79h3/5PFrCYwbdWhi3MAmnBk3pILdrHkh2JU4Ci6RwSpOzitl6rDBCGjQH
Druck0AIWGZl4ecz8EDh01CHQTIXeQBVUMHJ85LRvF8Q6rlJTmcpjBmbTV/WINxmy8114iLD65+e
SL5Sff1mbF8DUV2t3oGmIZmoNaBe9dmYZkZ25iz8rW+5ylvmAyl+TNHWUEfaiOd58vclu4d0/eJb
nVpE+p8dTMpmMWc8tI14EejevGQtL8jyVZOIz2eIDtTY/vPmaHTr9KTmm54pQ5rGg6Lb5yM+GD+F
qn+3tb5hxvNvhdUQB8vinNnNoemB8bGmJtz9HiwW1HWDtJFnYlfjkNe5JKMlIW/jbNr6mroZCaVH
56GCo194XkG8gQtsob4P4WyykeHcYS3HpaqOuAG3TgzytGyFKnTAHCxZ0Q6X9FQIVbGue5NFih+W
Lu6YxLeDWG38Y2DjFloSp3/sQRVku89MuPtifzuA1tK9KABLCsORrezpXH/R+2/h+8ZGoF9o0f0g
Avz5+jLIFfqFTAkt/J+GxcN8geDDd0h2XlLb/zrBhoXzwaTciFejOW71X14MtkAO3QU4W6kGLCQN
gh+bnCsunqKyjPjgTU6Rg1CqdjHI+1INsVTuUzudpiCzMlHiG907BMflWRJ3nghnRGQ+5eeICLLb
CCuzmh4rBCRJRARW04eZtfk6jYtb3W6u108iysx8ZURoA35YfiRSZSfy9B67sdspbNJnq5ooQvUs
4ai2XSQ+snyxntzSOmDByvoKQQG/RGkglN9qfP9xmuBTn0P5zUZUf1xtD/m48kyAYzZIeGKhBS0i
7c7kxrcR6aPwlL2fkp1uSZsEkg7bCGtqAMX1vcFjO0qtq2uSAl50wjhHyxr8Xws0KbIJT6Isp3rX
gyMt8jdJHWuOam4QCP0Wx4pJraLdTiPF7dO2RDHwExVigcRdV0xKUVAii/TboSDLmV8f8wg/PBue
VhsJy7Yv9CW7uj9WuCWLIzC1BTK/Yx61B3xSjn32uCdI9dw+yILDTau/thWMW1Xm7N+0/CXahjnN
NWSKHOAwkDCJX3Gi2mLH4m4nSoZ4/ZfAKqG3NDMb1a+yjEOcVgIrEDPN+pvYn02ykRqvtOUvapW1
UQ/BF9UC8m5/0VKfsLKJuz7sv28rt0IF81fbqXCe2bqbu4uk82ZVOcuz/oobhK/JVd0KzpWQ56ak
tyQ6s+w8INm/ZD6oh3wR38NaqyIuQqWAhf6fhb7BrZ+6jXNOWnMc2+PkdixwmZx9KWUBx+n6pHmj
a/djrLWXIKgfBxG931IQTDVD4G7SfVyyHQqG+Sn0JQRptmznk+2G2MilsR1XBn5sUi8KAw0rtkiW
ZQGT5U2EBdtNt+308ArqMkN5wedKE2Ugpwb2Yy604gMISlfOd3xFVcIJMD0kPiPYQkFirmHvSQLR
tyULaC4OQy1ef4dMDuGOxWnux5Wlk+YFFyd5E3yTGIrPR7wCqnigKcJqaubvhSsycau1Cj64Qy7U
q7DTzNEAIfWUH++A1M3PbQ5QnA0JbxK8sQ3QDoEfNivbWmdvdFNJ/a80U6aWvd0iI90wqRz8jFxA
vqx0uMHkNlXuulZ39bRWWjo1xS5i6wsZB/9wuuQ7UrRyLAx7jqKvYDwnd4S2Ab1ASaC6CAJmCZzh
IAMNwxSHe8NFagss9Vi7sy+d33nupEuPhtC+mtdUz2OXRJgHC9Nex2c204yJzE1+J2G6StuYar21
OQ6jUhVt3O/TaGBFITvdE8cJlwocnfseNyNFzh8NYC1CXf2Rvh8B2/7pIrjVgMqAB4D8QGkTB+Kd
o55ka1bfrrjrJv2yHM86anTs5/1b46CQ3Q8b83/xK7QJoGiCS/E+DdCK2Wxd+hAioBGsKe/9kAgv
jcYeG0D9zHXjddx95ev8picBec1iZLEIchYEpnnilKYopW6dGNSi1143DUtQrrp/wFaFqx+YqmMw
OtlmVxtQ9MBwAjfGW1o9hSQTk95BD/R1i6aZbe0ALacqEoU3YvekOfb+qFqEj3MHzUtRVIIL5H+K
C4gpn0bX/EXes+KDrdkVMu2OUqPUj8S/59TYcfaCnBwu9OZM4qA97BOZwh/fcZx+jw3wvh6esFYv
eGQsvayojTQST1wRXb3JZtbK242vRrncEifK2GdUoAc+leE6vfNvhcV0QYFQFxJFubHscGuTY/ic
5Apj0Ld4EBsFaX7HYqhkhmfxrDg7IWsHIEiLCpiKalpjvcnbBpSH91hQgVdM8h/suakeSBA78Nrw
p3uAWnHRpTV1050KmZDu69khd583PUHAKi947g7aFCDTDsAZ/XZAFyEcxCM2eEGJddxgRopVSJNh
Sju8jMBRHzXs/vCTBlqKm2t6jBK+8Gur0pclnYaFYtll7zBbCR09mwtukokzJ/g1p4BOGW7inXZU
groU3jZBy+tetrXZziSqUKx1eVTK4BpPey4mFecLaprQdKJ4sC+Qf/EB1akhMkELOlgB7I/2pOhS
5bwyMR+gD0NYOW7bielZ5DZyrNZMItgEuo5TCG+C/xG2Xbwa701raPbXN6JnL1CcnKq8Y1QJ+zOM
daFDsrOeQcZd4IRu1ancoHCHWrrR195JSILESW5eL89PKVf0Ux512puFaLVfFlJuo+oJFyiRbhJj
V9TvVOF9QbOiUKpNFUEO+cPsDoPgvgjYd1a3T3Avrk2oNCOSV3lsZV9O8Vs1BCuMcUbRsG1CnRi0
zOtINmyUyZms1BNzI/rIO+Flvyj1bN2UiaOoKPDs1n/kmCxAXnBHJT9R447MSShW1/fz5LR8eKaW
3qj1WXDCtZfimJcdyxPjsVTctguIP0xrO/mcnZ4dw+UznTwKmF2MIVM+ZRkxGEWr3Vbw/kCC3Msv
VOv+XMurJph7NMADukVfF0zjeY1bbBnxuAREpuNe+4qTbwZdld8a9Qnj7KhwiYs4S/gRzMHijV2K
PO8D7/piNiIG/3LoT/Mpz2RE+B+evpu968goUdYBbC9dr8RqTzYl+wbnjYESC6WHmmlsAt0vAYwR
VC6dcFUjB8LVHTW1iK0NKqQ6X+Rn4UUu9VWvxH674MPQZxh4DP0UdvOfXvcIqR6iK8UPKIEzqboI
J9SL05bgxAff28UFsCSBe7PRNjI1O6ATZIF1xop0Rqw7Pj+RfFJtAEUODSCIbWtdYJ3Ny9oNyU/m
4tOvG0J+zU7zdda52WHKmL/QIPXq73rjp0ZqCkGfFjTAdLZt3NvV9TxepZ7AUH3/4jzxnUy0RNPi
WP40UD3w/2n+gIOLrFHwkcl20CANrUBpsKg0ZzX5mBtuUS6/Z5fePURV/EhiFH2LcEM6SLVm6KKD
TYNFLr2nGnTLGpGTu3qIm4iwv7eJ8b0VUGj8wlr/F6PvSHt0zy/ESXdHMmZJAei2nYEXjOyLca9i
ej/XrAjIYOwhEDn+tWtLq5C1yuLeYZlfaDIcNpN+MuSluMXOBsDgbotGxqRfTcp77b1rxpXeOtI1
DYoW0hWRvhyDU5HwatsP86sPvPwGNg9r5AdGfC4pjzabYelhEa8vxt6vr+kNQaAy6Sb6bITFmoen
KdR0ffDSlkkJ4BVmKUvpf3ZHNddaBxjfqLRVR0j4kLj/73xd2c6xeqlHe3Zk9s0+kF/MLQkbaV/l
qAyjS0jbR73CwzTQEPqKNJvh92r+rbl+kshntzA8h8jmItqVweOadbHcMuUJGgKylOkerCjONmF2
RjdpKU5LSG6WBsdZpg2+REgMjIg21KD5oWH7EDlG5xlGjtRtMDXvHNoA8zECARTIAFJ4VDdGAgwQ
pV7JadUAGFVItyUSjYV0ewHNxXZyHWy05/3nUwo62ljecDa+c8ND9jcCgSrzccNeUI8pdR9nauT5
/OLVbYbxBBSmgOia7i7g+VlYIwrXHzTeFkLazhiz2nCayeKZXtK3+7Bnfvl+yzKYMKKa7mgr8ZOv
pCWrpUcoxWeoAUZUrcye/JLJeMcumf98hnU5BsvZPZrqyX2zA61Pr5i7kZsy9zSQYL5VHUgM5fQm
NlPKeplKlAqkLQ3Wyn41HIdGvUb0S3mJkOOF8/2ZeX9gTd8wXYhoX+P5NSlOKPwmXHOCYmZM8Dsm
BbaaAyunCz3FJeBiUNyJh5aRKAYvyPR2EJVC2Qs7aC0GOCsjIlH+JpNq/z8M/vGGnj+nX76tWZVI
dtUVa0hhGsDdE4/wRMRskvz63K0rmRJLUN5zCvjeWqpWYv1/S557UMiq0sT5Vr0YsU9Qso2HWXpz
Z3WMFXiYocOqpuDR9CQJ0Kw4trngwJZwCcx/Omq1Alk59QibVW9yhq2ueu7/7xP/0HK4eWb0Ojce
r/mliiDXajbZ7+V+w9uSPx1pskvjb+DmGAp7u8Jk6OkBjXn807iGZTmbKjjq7SHwWRuvHfPFOfGU
5/h9r9JkKVzMRtYAlaj4WD7dokqYz+CQ2XxxiWDXBxVQ4YpsMVp3UAC1d15DdkULj3m4wmjMcZl4
PFExqAettEN4UtFCYJ46FgKRVwiy1GvEvSFHp8CJ1ZrOO6YXNFBjd2/QGTJ4AE1arOsnqr6rhHgX
gvDqEUboJX1w0Y9r3QeKoj4N0maP9FDOtOZ3LX7c71dBSP8rm0x+1YYaDafOYSwPrHELO2a/Zz3f
9cDUtQ/TDnwcglj00Ua2xBf4iG+xFC6Ia+ERia8sP4p45ae1pb6RWFDmI1Z7TzzwGgx/INHgE+f2
hA/OSETokUWBl9slQW+/1WQQ7aE7jDJcK23uBtrJIfUEhb6zPSFdjkvtxo6Jgvf3Cr8vPuplniCl
m+TCiQL38QHBGj/rWsrAC/gF5Mp31GFey+B02a4Lvg+6+ZvF/zk3ue8zTRjm3yJGSdALoqLo9NB6
z7QlWGRYkIF6lcaMios4HFt8nXEG1RJ/4/rdkQShHQfxqI2Q13Vsq3ilV8lCD/gQ6ZOzeUoG0qpD
XD/G3wtf2LVk9pcl/RqC8tshR9imKvqgVd6zfTumVBoG8ip2w8bg2A428tfpZ2y/9gMxJe168GQr
0LNWChjd0SsT4g/kGN4LYCFIy1nx0h9G5U2vmwF89vhYRKdgSDCLGE5vyF10NlhvZaPv/mJusDmq
eH5NyQ/yL75lkjBl8wasiRd7rFaMpF+BuzaJp/zuG44JQtC6QjHiAoDeuac5pRVsB3ckJbv1TItP
+QclLLLJLuNOgEpc6w1aCyE4IiAWN6m6HPuxbl//p9/BdXKTrql6tCl/f3Q2TWSr44DvmkmjZ1+3
CFfbhP8iiMbm9nL+iPKLkWPBaHPgqEr5HqS5fdSbmU8TvueJMCnq1tTBXG1Sbul6FVDoP4RsU2vq
heAq2fixZAu8Y8JNmuuYkJR8KMm6LHGqagIgfuwz9qpQ0B5Rv9RCaE2UDE+aM4xeMk17fZcl/4qt
AW4DH9mgNSwBUcr2L7Bt4bP8lZlQPu+FSgGU+9EJvHOx/P5GGgzy4bMver8CXSU2OJJYpOf5HR0h
EfU8LEAja+IE2Op5u3GCljTHg6jRJgEUYT6SvKIJybfCSZmOAvu89nw+gb9cmWZ8Zx2jXuoqA5AN
JtKlT2VtwRAsUSV9EzixqUDK7Sf9Zqq14NiNOC1JElD1ZooiDvZZGRgmr6Xm2qxa+bcRRmegnDCT
gH6GFM4R8CLKDRFKig+6YhT1DT91BvNbBXqn20cEFhWPF6NNrw7cItWjOVaLyqZWSIeYps/qVdIv
hmB3mvqv4+iVSAcalGTxsOrpkT3oUFp1xXAq/d1sDqUVBQv4hMqtCUe6RUzWR0RnPrPYqPCPLCcW
LntkeeuFV1pI3LGIOb+xFM9hwukw4eZ91Jl2CkNZaG71J41mHrBhzdxcHwxu8VJF7WsGyXj775MI
EG98pWUkfvco3yfq85mn4iTT+aXx1KhT7pgWkcPHFu7kCEx0rBhk5GIUKVe2UJhz6KYPWNq80OwI
ujEOna7lH2aNg4FCQbjcvTf/26G+o7tUWuSQC3v0y26G9xDlxE/9dBWbd8HMpRatb5bSrhcvrzn8
boN0VL+0UYfXhT/8fzPs0qE/5rnxDvQJF8XL0xwv+8F+HKDZ2vF9Ghff1gphGyJVh36xmcv4H1jy
7QvvqSgQdLZLa6u1WbOT4cmgQwjvJWwr0Uln5jQls0Cn2Gk+3MCAOEsDA8+zoyj+4yZUaiz4AHjj
I2/abjIdqyHqtkGNiw/k+q1PpXdND9zHpEaTy10GVGlbCi5M+LeqDPe+d+JhjZKgLo+gAFTdqSTf
g1vWF5pfXrFgw76VnMW5qiOP/YONUYm9hcAzAMCi8RRsIWwG2SkIN7k2qfDecYLUUD/Ut3ONT8Fo
XebeKDAzN3tv/S+bkjECzKmKzLf28v0ttfYwzDFLVrQFMwSzAgSE+nak12EthxPAJrYSvRj00HSO
LegKizTBm/UsGLFlMTsPaRq5IUh4j/gC9R/Tw0/u7ICPhw/mXxTBZqqKAH0KlIl7UkhUTrTdvW5z
fAi2gAS6ngqh4almEkFe//0CEsO1kT1DBS3oclKw3jOnE4p86Nqf6jxG9MYLv5fiVr6SBPd5OTx5
Rnd+3YmRwD3crgETluajV9Fd4XtTvED9rlNFcI4Wtds7kTJaosdA0+CdKF6r98NdcURt44zry81x
q9Zn37M2/tN0IYoq7vbGjr4ZRTbmiBsWj/YuGfjRwig5YjFAqAx5zC6yiLuhTDqCwfcH8VoBq9QN
0LvHKAzlh1iQGkQKhtnY3E+Rgz9IVAsgtx9TLvmmgTj9JH8735nFe5ZybXZ1vonO2fc5c1XL+9dP
A+hWDUzP36aFR66Y7jxJkjxG38TOWbY2WN6vFsKZtHsrmj7duDgI6b5L1SPOm5LIVcElxHVOxcYu
b3C8J9iZLIbGXrGUnQ7J6EgEyIOEYPNluGgrtysHVGH8UEfEWecB23yubBJdp9VBUmxld5Huc5dj
uTQscI23A1k0L13MCzszNDwAqMCUj8NAGvSoSea5Cv/uCtK7j+48yRxVwFDlJdYG1UmcOakvQiNA
qngxecE8q3spjrYFi1HeNkUVqkzhfem6C2JjVS6yJOJr1EPdFbKbbDEGHD4Ig2w1M/Yl+RANuLar
Vuh9xMswVdbfE1kPJBDpkh7oYlWLQYQcERvqBumrGFy6WsWGAUHd5amXV1j7mt9UvOiMy7u0WFWT
GcqHacII0Wu3xu0qDLVX6J31mX9gNh7KoWSuSBAVYYaghBZnacIA42az0UAhhgsVHl1ZxrKMxm4t
Z4qgNEwiPq5deKRGF6bIZ1qkHfsY/5SfKDrwA8HBfvl+Vh0Lgtax4UoDo0HI7c4kWP8aYsvOaXnO
p6Wlai+tVDBUw7wpP1RJi7/mGKcpyfWwcAXaQK/9mDZm2EdYndjrbr1KVehAXtpKrkPDPok4JDgW
im63pfNgElSv+SktKIXJUeM3DHw1iEPTYqwbHI+Z9yJkqpGq4HMM/QYeNlCY+nChhZvbXD95CiSz
xC+Fy0Fz2rVnSV7cDk7q0kzUP0/oSY0AO9CRgESH6RJj+N8prlWfBoFilISwt08N8/9GazBS4Xsj
2zdSq9S25NxnYpdnQQUvOioKOEn1EvB23x1ZcwZU1xPgwpy3qFBzyWhiglebi/UQjyfcyTQCZ21u
ZbRKZub5QEIL/MAb/SWQ3qUxPucsnffuJKnpJQqURPpDsoG8+9+ccOdvjQmcYs8WlTMvHw7rnPXZ
9Y/pZYKJCGaKrBm05pRbTb8HHdpIlDV8nqaE5bJqSpvlEKnHrh5C78zuU8Zfk1BWvAFADldCfpsk
NsZ6KIDItBfsq27eq63L5hPGP32ujYQxTrSp2ChzOtaLMxkEqy9XgQIYtPDunLdEKgcI3GuaKsvh
thOj20oKB4EcBBMJd2z6G3Wiqvv6n/t354NJ/kGGSLqN1DXEf8NqprN/peYJ7j8CreenkfBhggNd
q2NS42MWHEX8qkLokmvIA5Zw0IYjlU4KfcdHmkr3MTq0OUE8Bh60eSzOvE9+ZkM01yL4DCDs7jF+
Le6uCGMqcTDYGccQ7yXPpYYgwvV+rJuf9Hgnbc7xlthfur1cQ1rvFDHhHXf1UCYfyNdHktEvntEn
WsrwbXS49jqmTG2K3wNOtQL+nBToOj5EUhEdgv91ghUAugg4bsFThYwwsmQVaFVu1hL+kRcjJ5a5
olROZIAaHrt5mZ3nXxapHHV0bmlxaQWmUfWgffXyqwkrkQ0P6FjJIPnCcxzayj+tJ+786haYHOVI
beEgDsJPhmj3O3AaH+1uZH7B+oDueCVjca9AOl4q6Q/4Zy07QddKgc696/3ph6yYsEf+ru1nSliE
lI08JVWHlkE24M89pZQuiIVfyWGqBr+v5Ijn3t0gs5lWWlP2el4PUOb38lMcCfDqZ0029RwvOQay
+48BkQ2E2UfY4+TdX8L0xhMHoK4zWd+2yaZmQN/He4S142ZSyubU+eqnnXmDJ/+yC6wD6Fbc7IiF
l98KHTyPy7fEMnQdsYuuWAMur/mMlnfERTxfV/TbXwQ39qjZH5Cs3Xt0NT8G3qUegM67ZlzkFi7T
UYxzfOPXt+R06cUY4uJykTTA/G4PwMSIkmI4UkHLRGoxMqtVF9pL+Kkk/wga32/CRCBdV8xRrZ3n
bnr1nB27xp92OCr/+cqapZAUVHpR9cKHoeW3VgbN/0DI4nifEeXnJOB7yd+ATJulMNnqIVtJvewq
eXaWoJ4Vp3bbgjv6iMkXkGOIizTaWgV9ok/0kyhoRNufZgDU1+QhvixhF6ijb5g8lnCj2p7gdNP6
Mrkd3xm4logyAWwa1qs6ooZD2nhzCa2hwlVc6zeMAFQI24FLSTG93kuf3emZ85EKnna9+YNIAQPM
DkcD5ORSJYjJoZ+FwYupffjgSshEfe591/pgycmd/ukUi1L1O9AnN3U2CQQuqnT5FV3ReU80q0V4
VWw2rS3GPq5fQAuhGeXv1HXVK3GdX+9fIgCarKXmImJOQ7ox4isGP8dXscjgI0xSdN3T5OTIWfK+
70hsebBF0LrBSlQajopu+v5tQO4rDpsCQa8N+xKac1ia8K5NCB6O6Eq6ZsqnngPljSvNnUiOu5CO
e3l4dijOeg9m7x0l4gPiuh07L3vnrLlTkHQuAIT3HTOnW4CP4KWGlqkcokqldxVwv2BgbB0EHNZH
d9uPLQfbSywbF0II43UiDIK3GxX0hpNvNlA8pHbmYp5yLBbi5Amt4ugi6wA+ctTTluBsBTD1EpfO
CE/Gjw/wq5wqSJaWphamK5AkGuFT5E6Q6Z8fLUihnyqf15Nni5Eex7vRI9n1mkK/09c0+JgzgATG
vQEoSbRSvfehzL16Zi/OrCS0VFKjjbaOMCfwJRphX4THw3iM9pD11JhDoVNebb2dO+nntnRWnBlb
9SSzHPMJG3J19CbF/PMm4xKeVpBhZWsXERYcANCTCFyHasAVt/kjbYfMWvTHmrviyzAWLo0hOBHH
kxa9zFAmYAa7MXqrD4yNszAhIylwwzDlgHL/x7D8zSBV9P1JExXP4SjiGp4dc6aF0mVsT+Fq3y1G
73Fp8LqSmdwn9lQuy2dEWAVQTnDFZj53Mg7NPYObMphKfD9BGA3+eCRT4t0HjUMi+RvLNHAREX3V
7QhsKTh/polPjFAliIHrO9Puhz+uxi0DGmimEHPGZJZhXBpMS31tb8NZ0CK0nLkd1LM02AQy1aRY
RRdXeXviBkEb2k6jeHlk9/pUqD1b1ilMIhzpwAUu5AgIeEg63LHPz1bKlCuOZSpXa9dcSMW9dgKl
tBoYMBOCKWfBjhK/4H9akAv9EDaxP8+uWfmZmnROnHAWV3cLIQ1MkEwzVO9ZsxQO53xs3mXMaKUw
aK/N5CwXrzt/pDnIC+zQAMsA53YqMMnHz2zDOA0zB1VyQx/4+aJ+2R3M5DU48/Qu1LPa/ChQ9AdL
DKJJOP0GVxO7yY8Nadsz8SJrNvV+ctKQ57U6JFHktMT11A6k+SWyFK4uu2np3rzzpEOxA7e2t6k/
3EKox02Ig6+TtWBEK+2VnOezsfyyb8pP5DGzjtoeRl6hICOwv2FlITVATFV7ojXBmyIe2zm9eeoF
2SSO0mW+oKJpqxYRODa/RukEafIutqS51bP2rw3aHOx1MBoF634/8NsOiZwuWHi6J3QH66aKK0mB
yPY9yU9M2tGbiO5ExCVCCw+SnwgJXShFWd4/5Ej1ZvY966Ffm151iDaXn+g9NVMES+UqnNGFpdem
dwv2Nr7xGRbVEEjlWMYo2Bps5BZ5jIW7atqvSHuTDNaKRjHZqRYYYEkbx9dxQDl97bf9W/u7FSM9
NZZlKBy+706J3QhjlxTsi9VEWP/QcDgOxf2VT2zRS+nCsY1XJmwdvA9G02HlPhcmgty6B4/Npq14
q9xXvcvm8R0BMRspzsqrkcQJO2lNlimyydJnLGRBAZoaEb++QpiKR/qkh4ihCBl7bhbwelpDYJP4
o29mBIjiUoPwpopLTyel9Qc5RirzgLCfMXsunhSF4cv2oiMSprePu6mshxxRaaSieLARBjH8tYHa
yUrpkUQNXgwkex9MPw4u8IUoQUeLmugzOhvUQO9aJVpyaFg1cNwYB4hXd2/r2UQIxtozebm6eFuc
IfkiTvJgJ0dwUZjrOCx2fmxAS9WkpsgrIvyr7ecPR4OFP1BazZ/KAjBIz26gCn+PuXLBUnrwXVhW
9U3fvWxLSGMVLoCiraS6eCP4VWvcWCLffQ1K+ZyV3gNz/VIQjwAnqbEdzJgUgmyeDejGFonb30Lo
5IevDve9AuDJZ5qsp+hWnGcmWV4JCIqCrX025/+B5b6exX+0y2lh1ifI9O20Q/9Dqy3wLzJOYj1V
BeGgxtUpE9q5O7JVVOiC8LwncyJ4jbBcw6cbtWFTTX9jV48Qc6k9DuXwCi8EM5RzMGWEUXqhYzFX
BFDacvdLb8WQrhmWgnp98xZwh94UuqYhk8jKOxdGYRR6p9VwL7NiJm90OzHwy5ZrUZWIsoDItZuT
vRZmYWl1Td0D+4cZUQm3U8fEe4YrTytjuLDTbovamHav9+CqWlJ6YQhwwEE03FBdwXFHgunb/sEx
QfA5sJkoxzy7Pxm+RObU2UA3qSWg7rbJMauBIG4NSLq/A+pCPvHhaRxv2lx2nYy6tvRYWICBlum4
gYxKpNeD0sHZppbI8msgokTdXp5A4YFf5FslI8g2aPAmuRwrwJWhf0PjuS6E36EK4aZI24byD9Pr
XENjrnosAw+uKBppzFuBcZcYRHNxWgIkaA3rxWhN4XwAxqbThmEpJXAQiBj8+LE+31hk0rYg7WEt
Ic1kuiMoeTeA9O8U10ArzPxL4S3G/vlSaUQRilJwQ4+G9rxMEJuXHdxtpLDvf3kWbLQHxfrSX/UG
qoUCGps9wmd2bt+1z6fvbPVgLC06qGnWdKfIXpTzMO+kD4+I4GD6C2r55MfQj9sy3zeryGqoxRBv
MW2OISTpDZbiLrWI97A8IUN301QPf+qgjzk11M0kM0KMDChsdCGdFV2tw8TjxyNDJqBw1LS0KOhO
wKjxmRrmZTM8l2tzBbm98wLaj9IOV+4t8ymMYv81EdXu9bKosmUqo5ITVzGG0wtlogVw1TgKBBXA
H3NMjvVGh4s3y0s3kmMo40HFmuTpn6jkm8LLTPx6qECY2pmyGqX8uFoQAQIb6mx3/wzi32cFHJzt
aJrxQ0gKXGYcm+cO6xn2zTpoU9KW5eKZll/aup9V0zns0OwrO4FtBCMIht0uiGp6GLVB85LrxJVt
u//2Wo2saf1nXkB7Zv307pCdx6Uv7wPpYJaM/P0pn9Cp8HUw8Tbh8noUeSs8tkxLKgaWh0TOg0FO
GEgmAQ5WVb7xirmGsI+aOWyPKYhFrzestGsZFZq20+bDg23Zq97W0u7gsXsiIkEAQr0uXz0I7Dtf
k+kRDg7djaF0+7LAPe7BwVp1heMznQDvbh26nNMpUVslyc+oYwphaBkdVTVHPPdtD2PS6vMNCHqz
S/z77G0iV/nklC/Z4a8agGAeruYJnC7zwd3nYUgxNIYvjcFlS1d/o0MqfnRBOW4QSHeZIrlEoMW+
cxJkJVDTE33s2l5qYFSVI+AvAXjOTy2N9LtA905n5Uh04gimqPiX8Ffkqpqy3jx2cYtqzqOHAtN+
9zXckJcLpykQh0pB/bJGIe54jlAgo7zAvs0lvCxwv3MPQrA+4guVXK7UW2sDKxBwA5rrRsvUlo0Y
737QucfPIv+zXurstRHBBaZmmbkDGq+eJZ97LwrdOX9gdlaTlb5IRGjD+aZfhONWIrryTG4s5jXd
tofx6GnNBC0sZpbj7/LwE8F1as5TcxujQ8CPjaJyZH67P3Nm50ZDhaD9fKwDhiAhu/GInZqMhkTZ
0CWhMMBAatVxqeeOGNIQclAOl5jUGrX9N55eREalVnsR4pJlJtj7LUz6PwK2iOhjIKiF0XOWWUtR
Wjj2XZ35ukYZVWp03R0bCHuEhvbWIeGLSN2CDn4FomKxgd+1lPF9HOZgsXZsxglv1jzMhVALtNsk
2LrCywrfQH6QJSVuXcog8SI98rr1hXFE4klnpfuq5nQTRfoJtJWYlps2nA522ArFfgdMHw9wENUd
e4Ua2VNAUohdNplTDxTsGmLsR405VKYOWY3cKKwJQGlUnqTSK7YwwEFt8nOw0meeoA1LYluPpsZR
4Ggk9aBBe4DbN1iqiKMxX2GdAoYfyIItAIPRYdzVKnGoQ4Yczhyvpc3TaOW4V98BDitpjJEZKWdU
CKGTFQAeujp4r4yJmWXeh6IuTfWiXRuCCX0ae/geegLkvRTeTZShVG0X7Lh9n+tW1uC5i4CDJu4M
lPabCDR9I3a5hflEkcVQPgtecIUg+yaprlShbxs1hhgf/g2ZE2yNdskqENtIf1KYvgvULuNj4T5H
IMQNtkxoDgPngY240tjEle+kHpaCCJaam/ncYy4CWi8tTiBZzYs/1IiHZHm6tsZGgoTJJ47RDjKg
7BUepuEC8x3qyGcj5qLb2L28M6cqTZwQxnGDl23lDpYuRVMvYDTSUK2XtVsq9DcSl6A1/Xt5WOjA
vlrOZeLCmatlJGGTr4XYYsEEyCIi8HpAhTrJkJM+Y6IoteXf/nC792nIcrY5nAs0A/p5+/EmbYBr
4Ht17ykTEBUJjAyaUJGA4m4HduZ/hTIjN1UZxkuq+vIfnaftSXVtlW4SG1ZIDwDmvJJ5vemQUGHB
7HHegrfuyx6rR4yyseXrfd6QrsqV9K5yVlpIWlrGM99HnYM0eqEetR6al1y687peRGODez+XO8ly
797vcYBTm0u7zoyZmrU4/gpDKfVSaoS42WvHeqclvo7fnUfOWzPbEoj41XBszT2WKZ7aFzVkIN07
0RiVGs1jLWmijOEyAIT74ktMlEUuFnL8
`protect end_protected
